magic
tech sky130A
magscale 1 2
timestamp 1739131682
<< nwell >>
rect 3359 1495 4732 2130
<< pwell >>
rect -928 587 4746 1434
<< psubdiff >>
rect -850 1333 -790 1367
rect 4618 1333 4678 1367
rect -850 1307 -816 1333
rect -850 699 -816 725
rect 4644 1307 4678 1333
rect 4644 699 4678 725
rect -850 665 -790 699
rect 4618 665 4678 699
<< nsubdiff >>
rect 3402 2049 3462 2083
rect 4626 2049 4686 2083
rect 3402 2023 3436 2049
rect 3402 1573 3436 1599
rect 4652 2023 4686 2049
rect 4652 1573 4686 1599
rect 3402 1539 3462 1573
rect 4626 1539 4686 1573
<< psubdiffcont >>
rect -790 1333 4618 1367
rect -850 725 -816 1307
rect 4644 725 4678 1307
rect -790 665 4618 699
<< nsubdiffcont >>
rect 3462 2049 4626 2083
rect 3402 1599 3436 2023
rect 4652 1599 4686 2023
rect 3462 1539 4626 1573
<< locali >>
rect 3292 2352 4734 2353
rect -504 2296 4734 2352
rect -504 2157 -374 2296
rect 4621 2157 4734 2296
rect -504 2083 4734 2157
rect -504 2049 3462 2083
rect 4626 2049 4734 2083
rect -504 2043 4734 2049
rect -504 2027 4735 2043
rect -504 1561 -426 2027
rect 186 1677 864 2027
rect 186 1561 264 1677
rect 779 1575 864 1677
rect 1485 2026 2258 2027
rect 2758 2026 3448 2027
rect 1485 1665 2162 2026
rect 1485 1575 1565 1665
rect -504 1495 265 1561
rect 775 1499 1565 1575
rect 2071 1573 2162 1665
rect 2759 2023 3448 2026
rect 2759 1665 3402 2023
rect 2759 1573 2855 1665
rect -502 1493 265 1495
rect 2071 1490 2855 1573
rect 3363 1599 3402 1665
rect 3436 1599 3448 2023
rect 3363 1578 3448 1599
rect 4631 2023 4735 2027
rect 4631 1599 4652 2023
rect 4686 1599 4735 2023
rect 4631 1578 4735 1599
rect 3363 1573 4735 1578
rect 3363 1539 3462 1573
rect 4626 1539 4735 1573
rect 3363 1501 4735 1539
rect 3365 1499 4735 1501
rect -897 1367 4725 1425
rect -897 1333 -790 1367
rect 4618 1333 4725 1367
rect -897 1307 4725 1333
rect -897 725 -850 1307
rect -816 1286 4644 1307
rect -816 791 -774 1286
rect 4602 791 4644 1286
rect -816 754 4644 791
rect -816 725 -804 754
rect -897 563 -804 725
rect 4603 725 4644 754
rect 4678 725 4725 1307
rect 4603 699 4725 725
rect 4618 665 4725 699
rect 4603 563 4725 665
rect -897 535 4725 563
<< viali >>
rect -374 2157 4621 2296
rect -804 699 4603 754
rect -804 665 -790 699
rect -790 665 4603 699
rect -804 563 4603 665
<< metal1 >>
rect 3306 2302 3364 2306
rect -386 2296 3279 2302
rect -386 2157 -374 2296
rect -386 2151 3279 2157
rect 4633 2151 4643 2302
rect 3306 2147 3364 2151
rect -386 1763 -376 1886
rect -324 1763 -314 1886
rect -267 1657 12 1943
rect 72 1710 82 1823
rect 134 1710 144 1823
rect 904 1763 914 1886
rect 966 1763 976 1886
rect 1031 1657 1310 1943
rect 1362 1710 1372 1823
rect 1424 1710 1434 1823
rect 2194 1763 2204 1886
rect 2256 1763 2266 1886
rect 2312 1657 2591 1943
rect 2652 1710 2662 1823
rect 2714 1710 2724 1823
rect 3484 1762 3494 1886
rect 3546 1762 3556 1886
rect 3622 1657 3901 1946
rect 3942 1710 3952 1833
rect 4004 1710 4014 1833
rect 4065 1763 4075 1886
rect 4127 1763 4137 1886
rect 4198 1657 4477 1945
rect 4523 1710 4533 1833
rect 4585 1710 4595 1833
rect -526 1611 4531 1657
rect -702 923 -692 983
rect -640 923 -630 983
rect -572 877 -505 1147
rect -442 1143 -372 1189
rect -444 923 -434 983
rect -382 923 -372 983
rect -442 833 -363 879
rect -314 877 -247 1147
rect -189 1143 -100 1189
rect -186 1099 -114 1143
rect -186 1039 -176 1099
rect -124 1039 -114 1099
rect -173 879 -127 913
rect -184 833 -115 879
rect -52 876 15 1146
rect 75 1143 145 1189
rect 72 923 82 983
rect 134 923 144 983
rect 75 833 143 879
rect 205 878 272 1148
rect 332 1144 401 1189
rect 330 1099 402 1144
rect 330 1039 340 1099
rect 392 1039 402 1099
rect 343 879 389 913
rect 333 833 401 879
rect 465 877 532 1147
rect 588 923 598 983
rect 650 923 660 983
rect 717 876 784 1146
rect 848 1143 917 1189
rect 846 923 856 983
rect 908 923 918 983
rect 848 833 916 879
rect 971 877 1038 1147
rect 1104 1143 1175 1189
rect 1104 1099 1176 1143
rect 1104 1039 1114 1099
rect 1166 1039 1176 1099
rect 1117 879 1163 912
rect 1106 833 1174 879
rect 1232 876 1299 1146
rect 1365 1143 1433 1189
rect 1362 923 1372 983
rect 1424 923 1434 983
rect 1362 833 1434 879
rect 1485 875 1552 1145
rect 1622 1143 1691 1189
rect 1620 1099 1692 1143
rect 1620 1039 1630 1099
rect 1682 1039 1692 1099
rect 1633 879 1679 912
rect 1622 833 1694 879
rect 1747 877 1814 1147
rect 1878 923 1888 983
rect 1940 923 1950 983
rect 2005 878 2072 1148
rect 2137 1143 2207 1189
rect 2136 923 2146 983
rect 2198 923 2208 983
rect 2138 833 2206 879
rect 2262 878 2329 1148
rect 2396 1144 2466 1189
rect 2394 1099 2466 1144
rect 2394 1039 2404 1099
rect 2456 1039 2466 1099
rect 2407 879 2453 916
rect 2396 833 2464 879
rect 2523 878 2590 1148
rect 2652 1143 2724 1189
rect 2652 923 2662 983
rect 2714 923 2724 983
rect 2655 833 2723 879
rect 2782 876 2849 1146
rect 2911 1145 2983 1189
rect 2910 1143 2983 1145
rect 2910 1099 2982 1143
rect 2910 1039 2920 1099
rect 2972 1039 2982 1099
rect 2923 879 2969 914
rect 2912 833 2980 879
rect 3032 877 3099 1147
rect 3168 923 3178 983
rect 3230 923 3240 983
rect 3292 877 3359 1147
rect 3429 1143 3496 1189
rect 3426 923 3436 983
rect 3488 923 3498 983
rect 3429 833 3495 879
rect 3554 876 3621 1146
rect 3687 1144 3754 1189
rect 3684 1099 3756 1144
rect 3684 1039 3694 1099
rect 3746 1039 3756 1099
rect 3697 879 3743 914
rect 3687 833 3753 879
rect 3814 876 3881 1146
rect 3945 1143 4012 1189
rect 3942 923 3952 983
rect 4004 923 4014 983
rect 3943 833 4013 879
rect 4073 876 4140 1146
rect 4202 1144 4269 1189
rect 4200 1099 4272 1144
rect 4200 1039 4210 1099
rect 4262 1039 4272 1099
rect 4213 879 4259 914
rect 4202 833 4269 879
rect 4340 877 4407 1147
rect 4458 1039 4468 1099
rect 4520 1039 4530 1099
rect 4458 923 4468 983
rect 4520 923 4530 983
rect -816 754 4615 760
rect -816 563 -804 754
rect 4603 563 4615 754
rect -816 557 4615 563
<< via1 >>
rect 3279 2296 4633 2302
rect -374 2157 4621 2296
rect 4621 2157 4633 2296
rect 3279 2151 4633 2157
rect -376 1763 -324 1886
rect 82 1710 134 1823
rect 914 1763 966 1886
rect 1372 1710 1424 1823
rect 2204 1763 2256 1886
rect 2662 1710 2714 1823
rect 3494 1762 3546 1886
rect 3952 1710 4004 1833
rect 4075 1763 4127 1886
rect 4533 1710 4585 1833
rect -692 923 -640 983
rect -434 923 -382 983
rect -176 1039 -124 1099
rect 82 923 134 983
rect 340 1039 392 1099
rect 598 923 650 983
rect 856 923 908 983
rect 1114 1039 1166 1099
rect 1372 923 1424 983
rect 1630 1039 1682 1099
rect 1888 923 1940 983
rect 2146 923 2198 983
rect 2404 1039 2456 1099
rect 2662 923 2714 983
rect 2920 1039 2972 1099
rect 3178 923 3230 983
rect 3436 923 3488 983
rect 3694 1039 3746 1099
rect 3952 923 4004 983
rect 4210 1039 4262 1099
rect 4468 1039 4520 1099
rect 4468 923 4520 983
rect -804 563 4603 754
<< metal2 >>
rect 3279 2306 4633 2312
rect -547 2302 4633 2306
rect -547 2296 3279 2302
rect -547 2157 -374 2296
rect -547 2151 3279 2157
rect -547 2147 4633 2151
rect -376 1886 -324 2147
rect 914 1886 966 2147
rect -376 1753 -324 1763
rect 82 1823 134 1833
rect 2204 1886 2256 2147
rect 3279 2141 4633 2147
rect 914 1753 966 1763
rect 1372 1823 1424 1833
rect 82 1109 134 1710
rect 3494 1886 3546 2141
rect 2204 1753 2256 1763
rect 2662 1823 2714 1833
rect 1372 1109 1424 1710
rect 4075 1886 4127 2141
rect 3494 1752 3546 1762
rect 3952 1833 4004 1842
rect 2662 1109 2714 1710
rect 4075 1753 4127 1763
rect 4533 1833 4585 1843
rect 3952 1109 4004 1710
rect 4533 1471 4585 1710
rect 4468 1422 4746 1471
rect -176 1099 392 1109
rect -124 1039 340 1099
rect -176 1029 392 1039
rect 1114 1099 1682 1109
rect 1166 1039 1630 1099
rect 1114 1029 1682 1039
rect 2404 1099 2972 1109
rect 2456 1039 2920 1099
rect 2404 1029 2972 1039
rect 3694 1099 4262 1109
rect 3746 1039 4210 1099
rect 3694 1029 4262 1039
rect 4468 1099 4520 1422
rect 4468 993 4520 1039
rect -928 983 -640 993
rect -928 923 -692 983
rect -928 913 -640 923
rect -434 983 650 993
rect -382 923 82 983
rect 134 923 598 983
rect -434 913 650 923
rect 856 983 1940 993
rect 908 923 1372 983
rect 1424 923 1888 983
rect 856 913 1940 923
rect 2146 983 3230 993
rect 2198 923 2662 983
rect 2714 923 3178 983
rect 2146 913 3230 923
rect 3436 983 4520 993
rect 3488 923 3952 983
rect 4004 923 4468 983
rect 3436 913 4520 923
rect -897 754 4603 764
rect -897 563 -804 754
rect -897 553 4603 563
use sky130_fd_pr__nfet_01v8_lvt_LH3874  sky130_fd_pr__nfet_01v8_lvt_LH3874_0
timestamp 1738199432
transform 1 0 4365 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__pfet_01v8_lvt_Q4S9T2  sky130_fd_pr__pfet_01v8_lvt_Q4S9T2_0
timestamp 1738897390
transform 1 0 2459 0 1 1798
box -396 -319 396 319
use sky130_fd_pr__pfet_01v8_lvt_Q4S9T2  sky130_fd_pr__pfet_01v8_lvt_Q4S9T2_1
timestamp 1738897390
transform 1 0 -121 0 1 1798
box -396 -319 396 319
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM1
timestamp 1738199432
transform 1 0 -21 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM2
timestamp 1738199432
transform 1 0 237 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM3
timestamp 1738199432
transform 1 0 495 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM4
timestamp 1738199432
transform 1 0 -537 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM5
timestamp 1738199432
transform 1 0 -279 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM6
timestamp 1738199432
transform 1 0 753 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM7
timestamp 1738199432
transform 1 0 1011 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM8
timestamp 1738199432
transform 1 0 1269 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM9
timestamp 1738199432
transform 1 0 1527 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__pfet_01v8_lvt_Q4S9T2  XM11
timestamp 1738897390
transform 1 0 1169 0 1 1798
box -396 -319 396 319
use sky130_fd_pr__pfet_01v8_lvt_L4HHUA  XM12
timestamp 1738899194
transform 1 0 4330 0 1 1798
box -294 -200 294 200
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM13
timestamp 1738199432
transform 1 0 1785 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM15
timestamp 1738199432
transform 1 0 2301 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM16
timestamp 1738199432
transform 1 0 2043 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__pfet_01v8_lvt_QCP9T2  XM17
timestamp 1738899194
transform 1 0 3749 0 1 1798
box -294 -200 294 200
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM18
timestamp 1738199432
transform 1 0 3591 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM19
timestamp 1738199432
transform 1 0 3333 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM20
timestamp 1738199432
transform 1 0 2559 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM21
timestamp 1738199432
transform 1 0 2817 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM22
timestamp 1738199432
transform 1 0 3075 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM23
timestamp 1738199432
transform 1 0 3849 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM24
timestamp 1738199432
transform 1 0 4107 0 1 1011
box -158 -188 158 188
<< labels >>
rlabel metal2 -422 2228 -422 2228 3 vcc
port 1 e
rlabel metal2 -896 637 -896 637 3 vss
port 2 e
rlabel metal2 -927 957 -927 957 3 vref0
port 4 e
rlabel metal1 -494 1637 -494 1637 3 vr
port 5 e
rlabel metal2 4745 1447 4745 1447 7 vref
port 3 w
<< end >>
