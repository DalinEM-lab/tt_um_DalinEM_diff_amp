magic
tech sky130A
magscale 1 2
timestamp 1738875365
<< nwell >>
rect 3404 1459 4739 2338
<< pwell >>
rect -928 587 4746 1434
<< psubdiff >>
rect -850 1333 -790 1367
rect 4618 1333 4678 1367
rect -850 1307 -816 1333
rect -850 699 -816 725
rect 4644 1307 4678 1333
rect 4644 699 4678 725
rect -850 665 -790 699
rect 4618 665 4678 699
<< nsubdiff >>
rect 3472 2260 3532 2294
rect 4598 2260 4658 2294
rect 3472 2206 3506 2260
rect 3472 1556 3506 1582
rect 4624 2206 4658 2260
rect 4624 1556 4658 1582
rect 3472 1522 3532 1556
rect 4598 1522 4658 1556
<< psubdiffcont >>
rect -790 1333 4618 1367
rect -850 725 -816 1307
rect 4644 725 4678 1307
rect -790 665 4618 699
<< nsubdiffcont >>
rect 3532 2260 4598 2294
rect 3472 1582 3506 2206
rect 4624 1582 4658 2206
rect 3532 1522 4598 1556
<< locali >>
rect -423 2296 4741 2352
rect -423 2157 -374 2296
rect -423 2027 3472 2157
rect -423 1576 -329 2027
rect 177 1576 278 2027
rect -423 1479 278 1576
rect 852 1573 968 2027
rect 1465 1573 1572 2027
rect 852 1476 1572 1573
rect 2165 1577 2258 2027
rect 2758 1577 2865 2027
rect 3364 2023 3472 2027
rect 2165 1480 2865 1577
rect 3404 1582 3472 2023
rect 3506 2023 4624 2157
rect 3506 1582 3530 2023
rect 3404 1572 3530 1582
rect 4598 1582 4624 2023
rect 4658 1582 4741 2296
rect 4598 1572 4741 1582
rect 3404 1563 4741 1572
rect 3404 1556 4740 1563
rect 3404 1522 3532 1556
rect 4598 1522 4740 1556
rect 3404 1459 4740 1522
rect -897 1367 4725 1425
rect -897 1333 -790 1367
rect 4618 1333 4725 1367
rect -897 1307 4725 1333
rect -897 725 -850 1307
rect -816 1286 4644 1307
rect -816 791 -774 1286
rect 4602 791 4644 1286
rect -816 754 4644 791
rect -816 725 -804 754
rect -897 563 -804 725
rect 4603 725 4644 754
rect 4678 725 4725 1307
rect 4603 699 4725 725
rect 4618 665 4725 699
rect 4603 563 4725 665
rect -897 535 4725 563
<< viali >>
rect -374 2294 4658 2296
rect -374 2260 3532 2294
rect 3532 2260 4598 2294
rect 4598 2260 4658 2294
rect -374 2206 4658 2260
rect -374 2157 3472 2206
rect 3472 2157 3506 2206
rect 3506 2157 4624 2206
rect 4624 2157 4658 2206
rect -804 699 4603 754
rect -804 665 -790 699
rect -790 665 4603 699
rect -804 563 4603 665
<< metal1 >>
rect -386 2296 4670 2302
rect -386 2157 -374 2296
rect 4658 2157 4670 2296
rect -386 2151 4670 2157
rect -306 1826 -296 1886
rect -244 1826 -234 1886
rect -164 1657 11 1943
rect 984 1816 994 1886
rect 1046 1816 1056 1886
rect 72 1710 82 1770
rect 134 1710 144 1770
rect 1132 1657 1307 1944
rect 2274 1816 2284 1886
rect 2336 1816 2346 1886
rect 1362 1710 1372 1780
rect 1424 1710 1434 1780
rect 2429 1657 2604 1945
rect 3564 1816 3574 1886
rect 3626 1816 3636 1886
rect 2652 1710 2662 1780
rect 2714 1710 2724 1780
rect 3711 1657 3886 1945
rect 4269 1939 4272 1985
rect 4200 1816 4210 1886
rect 4262 1816 4272 1886
rect 3942 1710 3952 1780
rect 4004 1710 4014 1780
rect -495 1611 4271 1657
rect 4304 1653 4418 1985
rect 4458 1939 4461 1950
rect 4458 1902 4530 1910
rect 4458 1710 4468 1902
rect 4520 1710 4530 1902
rect -702 923 -692 983
rect -640 923 -630 983
rect -572 877 -505 1147
rect -442 1143 -372 1189
rect -444 923 -434 983
rect -382 923 -372 983
rect -442 833 -363 879
rect -314 877 -247 1147
rect -189 1143 -100 1189
rect -186 1099 -114 1143
rect -186 1039 -176 1099
rect -124 1039 -114 1099
rect -173 879 -127 913
rect -184 833 -115 879
rect -52 876 15 1146
rect 75 1143 145 1189
rect 72 923 82 983
rect 134 923 144 983
rect 75 833 143 879
rect 205 878 272 1148
rect 332 1144 401 1189
rect 330 1099 402 1144
rect 330 1039 340 1099
rect 392 1039 402 1099
rect 343 879 389 913
rect 333 833 401 879
rect 465 877 532 1147
rect 588 923 598 983
rect 650 923 660 983
rect 717 876 784 1146
rect 848 1143 917 1189
rect 846 923 856 983
rect 908 923 918 983
rect 848 833 916 879
rect 971 877 1038 1147
rect 1104 1143 1175 1189
rect 1104 1099 1176 1143
rect 1104 1039 1114 1099
rect 1166 1039 1176 1099
rect 1117 879 1163 912
rect 1106 833 1174 879
rect 1232 876 1299 1146
rect 1365 1143 1433 1189
rect 1362 923 1372 983
rect 1424 923 1434 983
rect 1362 833 1434 879
rect 1485 875 1552 1145
rect 1622 1143 1691 1189
rect 1620 1099 1692 1143
rect 1620 1039 1630 1099
rect 1682 1039 1692 1099
rect 1633 879 1679 912
rect 1622 833 1694 879
rect 1747 877 1814 1147
rect 1878 923 1888 983
rect 1940 923 1950 983
rect 2005 878 2072 1148
rect 2137 1143 2207 1189
rect 2136 923 2146 983
rect 2198 923 2208 983
rect 2138 833 2206 879
rect 2262 878 2329 1148
rect 2396 1144 2466 1189
rect 2394 1099 2466 1144
rect 2394 1039 2404 1099
rect 2456 1039 2466 1099
rect 2407 879 2453 916
rect 2396 833 2464 879
rect 2523 878 2590 1148
rect 2652 1143 2724 1189
rect 2652 923 2662 983
rect 2714 923 2724 983
rect 2655 833 2723 879
rect 2782 876 2849 1146
rect 2911 1145 2983 1189
rect 2910 1143 2983 1145
rect 2910 1099 2982 1143
rect 2910 1039 2920 1099
rect 2972 1039 2982 1099
rect 2923 879 2969 914
rect 2912 833 2980 879
rect 3032 877 3099 1147
rect 3168 923 3178 983
rect 3230 923 3240 983
rect 3292 877 3359 1147
rect 3429 1143 3496 1189
rect 3426 923 3436 983
rect 3488 923 3498 983
rect 3429 833 3495 879
rect 3554 876 3621 1146
rect 3687 1144 3754 1189
rect 3684 1099 3756 1144
rect 3684 1039 3694 1099
rect 3746 1039 3756 1099
rect 3697 879 3743 914
rect 3687 833 3753 879
rect 3814 876 3881 1146
rect 3945 1143 4012 1189
rect 3942 923 3952 983
rect 4004 923 4014 983
rect 3943 833 4013 879
rect 4073 876 4140 1146
rect 4202 1144 4269 1189
rect 4200 1099 4272 1144
rect 4200 1039 4210 1099
rect 4262 1039 4272 1099
rect 4213 879 4259 914
rect 4202 833 4269 879
rect 4340 877 4407 1147
rect 4458 1039 4468 1099
rect 4520 1039 4530 1099
rect 4458 923 4468 983
rect 4520 923 4530 983
rect -816 754 4615 760
rect -816 563 -804 754
rect 4603 563 4615 754
rect -816 557 4615 563
<< via1 >>
rect -374 2157 4658 2296
rect -296 1826 -244 1886
rect 994 1816 1046 1886
rect 82 1710 134 1770
rect 2284 1816 2336 1886
rect 1372 1710 1424 1780
rect 3574 1816 3626 1886
rect 2662 1710 2714 1780
rect 4210 1816 4262 1886
rect 3952 1710 4004 1780
rect 4468 1710 4520 1902
rect -692 923 -640 983
rect -434 923 -382 983
rect -176 1039 -124 1099
rect 82 923 134 983
rect 340 1039 392 1099
rect 598 923 650 983
rect 856 923 908 983
rect 1114 1039 1166 1099
rect 1372 923 1424 983
rect 1630 1039 1682 1099
rect 1888 923 1940 983
rect 2146 923 2198 983
rect 2404 1039 2456 1099
rect 2662 923 2714 983
rect 2920 1039 2972 1099
rect 3178 923 3230 983
rect 3436 923 3488 983
rect 3694 1039 3746 1099
rect 3952 923 4004 983
rect 4210 1039 4262 1099
rect 4468 1039 4520 1099
rect 4468 923 4520 983
rect -804 563 4603 754
<< metal2 >>
rect -423 2296 4658 2306
rect -423 2157 -374 2296
rect -423 2147 4658 2157
rect -296 1886 -244 2147
rect -296 1816 -244 1826
rect 994 1886 1046 2147
rect 994 1806 1046 1816
rect 2284 1886 2336 2147
rect 2284 1806 2336 1816
rect 3574 1886 3626 2147
rect 3574 1806 3626 1816
rect 4210 1886 4262 2147
rect 4210 1806 4262 1816
rect 4468 1902 4520 1921
rect 1372 1780 1424 1790
rect 82 1770 134 1780
rect 82 1109 134 1710
rect 1372 1109 1424 1710
rect 2662 1780 2714 1790
rect 2662 1109 2714 1710
rect 3952 1780 4004 1790
rect 3952 1109 4004 1710
rect 4468 1474 4520 1710
rect 4468 1422 4746 1474
rect -176 1099 392 1109
rect -124 1039 340 1099
rect -176 1029 392 1039
rect 1114 1099 1682 1109
rect 1166 1039 1630 1099
rect 1114 1029 1682 1039
rect 2404 1099 2972 1109
rect 2456 1039 2920 1099
rect 2404 1029 2972 1039
rect 3694 1099 4262 1109
rect 3746 1039 4210 1099
rect 3694 1029 4262 1039
rect 4468 1099 4520 1422
rect 4468 993 4520 1039
rect -928 983 -640 993
rect -928 923 -692 983
rect -928 913 -640 923
rect -434 983 650 993
rect -382 923 82 983
rect 134 923 598 983
rect -434 913 650 923
rect 856 983 1940 993
rect 908 923 1372 983
rect 1424 923 1888 983
rect 856 913 1940 923
rect 2146 983 3230 993
rect 2198 923 2662 983
rect 2714 923 3178 983
rect 2146 913 3230 923
rect 3436 983 4520 993
rect 3488 923 3952 983
rect 4004 923 4468 983
rect 3436 913 4520 923
rect -897 754 4603 764
rect -897 563 -804 754
rect -897 553 4603 563
use sky130_fd_pr__nfet_01v8_lvt_LH3874  sky130_fd_pr__nfet_01v8_lvt_LH3874_0
timestamp 1738199432
transform 1 0 4365 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__pfet_01v8_lvt_QPK3U4  sky130_fd_pr__pfet_01v8_lvt_QPK3U4_0
timestamp 1738725867
transform 1 0 2499 0 1 1798
box -356 -319 356 319
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM1
timestamp 1738199432
transform 1 0 -21 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM2
timestamp 1738199432
transform 1 0 237 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM3
timestamp 1738199432
transform 1 0 495 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM4
timestamp 1738199432
transform 1 0 -537 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM5
timestamp 1738199432
transform 1 0 -279 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM6
timestamp 1738199432
transform 1 0 753 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM7
timestamp 1738199432
transform 1 0 1011 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM8
timestamp 1738199432
transform 1 0 1269 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM9
timestamp 1738199432
transform 1 0 1527 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__pfet_01v8_lvt_QPK3U4  XM10
timestamp 1738725867
transform 1 0 -81 0 1 1798
box -356 -319 356 319
use sky130_fd_pr__pfet_01v8_lvt_QPK3U4  XM11
timestamp 1738725867
transform 1 0 1209 0 1 1798
box -356 -319 356 319
use sky130_fd_pr__pfet_01v8_lvt_QCPJZY  XM12
timestamp 1738726022
transform 1 0 4365 0 1 1798
box -194 -200 194 200
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM13
timestamp 1738199432
transform 1 0 1785 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM15
timestamp 1738199432
transform 1 0 2301 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM16
timestamp 1738199432
transform 1 0 2043 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__pfet_01v8_lvt_QXG3U4  XM17
timestamp 1738726022
transform 1 0 3789 0 1 1798
box -254 -200 254 200
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM18
timestamp 1738199432
transform 1 0 3591 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM19
timestamp 1738199432
transform 1 0 3333 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM20
timestamp 1738199432
transform 1 0 2559 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM21
timestamp 1738199432
transform 1 0 2817 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM22
timestamp 1738199432
transform 1 0 3075 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM23
timestamp 1738199432
transform 1 0 3849 0 1 1011
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_lvt_LH3874  XM24
timestamp 1738199432
transform 1 0 4107 0 1 1011
box -158 -188 158 188
<< labels >>
rlabel metal2 -422 2228 -422 2228 3 vcc
port 1 e
rlabel metal2 4745 1450 4745 1450 3 vref
port 3 e
rlabel metal2 -896 637 -896 637 3 vss
port 2 e
rlabel metal2 -927 957 -927 957 3 vref0
port 4 e
rlabel metal1 -494 1637 -494 1637 3 vr
port 5 e
<< end >>
