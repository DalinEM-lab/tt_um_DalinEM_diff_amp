magic
tech sky130A
magscale 1 2
timestamp 1741206017
<< nwell >>
rect 3680 3190 4498 4148
rect -820 484 4074 2918
<< pwell >>
rect 881 5486 2401 6536
rect 556 3053 2692 5338
rect 3160 5204 4564 5606
<< nmos >>
rect 1091 6040 2191 6340
rect 1091 5682 2191 5982
<< pmoslvt >>
rect 3876 3409 3946 3929
rect 4232 3409 4302 3929
rect -457 2006 543 2506
rect 601 2006 1601 2506
rect 1659 2006 2659 2506
rect 2717 2006 3717 2506
rect -457 844 543 1344
rect 601 844 1601 1344
rect 1659 844 2659 1344
rect 2717 844 3717 1344
<< nmoslvt >>
rect 728 4498 1128 5098
rect 1186 4498 1586 5098
rect 1644 4498 2044 5098
rect 2102 4498 2502 5098
rect 728 3291 1128 3891
rect 1186 3291 1586 3891
rect 1644 3291 2044 3891
rect 2102 3291 2502 3891
rect 3916 4414 3946 4614
rect 4272 4414 4302 4614
<< ndiff >>
rect 1091 6386 2191 6398
rect 1091 6352 1103 6386
rect 2179 6352 2191 6386
rect 1091 6340 2191 6352
rect 1091 6028 2191 6040
rect 1091 5994 1103 6028
rect 2179 5994 2191 6028
rect 1091 5982 2191 5994
rect 1091 5670 2191 5682
rect 1091 5636 1103 5670
rect 2179 5636 2191 5670
rect 1091 5624 2191 5636
rect 670 5086 728 5098
rect 670 4510 682 5086
rect 716 4510 728 5086
rect 670 4498 728 4510
rect 1128 5086 1186 5098
rect 1128 4510 1140 5086
rect 1174 4510 1186 5086
rect 1128 4498 1186 4510
rect 1586 5086 1644 5098
rect 1586 4510 1598 5086
rect 1632 4510 1644 5086
rect 1586 4498 1644 4510
rect 2044 5086 2102 5098
rect 2044 4510 2056 5086
rect 2090 4510 2102 5086
rect 2044 4498 2102 4510
rect 2502 5086 2560 5098
rect 2502 4510 2514 5086
rect 2548 4510 2560 5086
rect 2502 4498 2560 4510
rect 670 3879 728 3891
rect 670 3303 682 3879
rect 716 3303 728 3879
rect 670 3291 728 3303
rect 1128 3879 1186 3891
rect 1128 3303 1140 3879
rect 1174 3303 1186 3879
rect 1128 3291 1186 3303
rect 1586 3879 1644 3891
rect 1586 3303 1598 3879
rect 1632 3303 1644 3879
rect 1586 3291 1644 3303
rect 2044 3879 2102 3891
rect 2044 3303 2056 3879
rect 2090 3303 2102 3879
rect 2044 3291 2102 3303
rect 2502 3879 2560 3891
rect 2502 3303 2514 3879
rect 2548 3303 2560 3879
rect 2502 3291 2560 3303
rect 3858 4602 3916 4614
rect 3858 4426 3870 4602
rect 3904 4426 3916 4602
rect 3858 4414 3916 4426
rect 3946 4602 4004 4614
rect 3946 4426 3958 4602
rect 3992 4426 4004 4602
rect 3946 4414 4004 4426
rect 4214 4602 4272 4614
rect 4214 4426 4226 4602
rect 4260 4426 4272 4602
rect 4214 4414 4272 4426
rect 4302 4602 4360 4614
rect 4302 4426 4314 4602
rect 4348 4426 4360 4602
rect 4302 4414 4360 4426
<< pdiff >>
rect 3818 3917 3876 3929
rect 3818 3421 3830 3917
rect 3864 3421 3876 3917
rect 3818 3409 3876 3421
rect 3946 3917 4004 3929
rect 3946 3421 3958 3917
rect 3992 3421 4004 3917
rect 3946 3409 4004 3421
rect 4174 3917 4232 3929
rect 4174 3421 4186 3917
rect 4220 3421 4232 3917
rect 4174 3409 4232 3421
rect 4302 3917 4360 3929
rect 4302 3421 4314 3917
rect 4348 3421 4360 3917
rect 4302 3409 4360 3421
rect -515 2494 -457 2506
rect -515 2018 -503 2494
rect -469 2018 -457 2494
rect -515 2006 -457 2018
rect 543 2494 601 2506
rect 543 2018 555 2494
rect 589 2018 601 2494
rect 543 2006 601 2018
rect 1601 2494 1659 2506
rect 1601 2018 1613 2494
rect 1647 2018 1659 2494
rect 1601 2006 1659 2018
rect 2659 2494 2717 2506
rect 2659 2018 2671 2494
rect 2705 2018 2717 2494
rect 2659 2006 2717 2018
rect 3717 2494 3775 2506
rect 3717 2018 3729 2494
rect 3763 2018 3775 2494
rect 3717 2006 3775 2018
rect -515 1332 -457 1344
rect -515 856 -503 1332
rect -469 856 -457 1332
rect -515 844 -457 856
rect 543 1332 601 1344
rect 543 856 555 1332
rect 589 856 601 1332
rect 543 844 601 856
rect 1601 1332 1659 1344
rect 1601 856 1613 1332
rect 1647 856 1659 1332
rect 1601 844 1659 856
rect 2659 1332 2717 1344
rect 2659 856 2671 1332
rect 2705 856 2717 1332
rect 2659 844 2717 856
rect 3717 1332 3775 1344
rect 3717 856 3729 1332
rect 3763 856 3775 1332
rect 3717 844 3775 856
<< ndiffc >>
rect 1103 6352 2179 6386
rect 1103 5994 2179 6028
rect 1103 5636 2179 5670
rect 682 4510 716 5086
rect 1140 4510 1174 5086
rect 1598 4510 1632 5086
rect 2056 4510 2090 5086
rect 2514 4510 2548 5086
rect 682 3303 716 3879
rect 1140 3303 1174 3879
rect 1598 3303 1632 3879
rect 2056 3303 2090 3879
rect 2514 3303 2548 3879
rect 3870 4426 3904 4602
rect 3958 4426 3992 4602
rect 4226 4426 4260 4602
rect 4314 4426 4348 4602
<< pdiffc >>
rect 3830 3421 3864 3917
rect 3958 3421 3992 3917
rect 4186 3421 4220 3917
rect 4314 3421 4348 3917
rect -503 2018 -469 2494
rect 555 2018 589 2494
rect 1613 2018 1647 2494
rect 2671 2018 2705 2494
rect 3729 2018 3763 2494
rect -503 856 -469 1332
rect 555 856 589 1332
rect 1613 856 1647 1332
rect 2671 856 2705 1332
rect 3729 856 3763 1332
<< psubdiff >>
rect 917 6466 1013 6500
rect 2269 6466 2365 6500
rect 917 6404 951 6466
rect 2331 6404 2365 6466
rect 917 5556 951 5618
rect 2331 5556 2365 5618
rect 917 5522 1013 5556
rect 2269 5522 2365 5556
rect 3196 5536 3292 5570
rect 4432 5536 4528 5570
rect 3196 5474 3230 5536
rect 4494 5474 4528 5536
rect 572 5279 632 5313
rect 2614 5279 2674 5313
rect 572 5253 606 5279
rect 2640 5253 2674 5279
rect 572 3109 606 3135
rect 3196 5274 3230 5336
rect 4494 5274 4528 5336
rect 3196 5240 3292 5274
rect 4432 5240 4528 5274
rect 3748 4766 3808 4800
rect 4407 4766 4467 4800
rect 3748 4740 3782 4766
rect 4433 4740 4467 4766
rect 3748 4274 3782 4300
rect 4433 4274 4467 4300
rect 3748 4240 3808 4274
rect 4407 4240 4467 4274
rect 2640 3109 2674 3135
rect 572 3075 632 3109
rect 2614 3075 2674 3109
<< nsubdiff >>
rect 3716 4078 3812 4112
rect 4010 4078 4168 4112
rect 4366 4078 4462 4112
rect 3716 4016 3750 4078
rect 4072 4016 4106 4078
rect 3716 3260 3750 3322
rect 4428 4016 4462 4078
rect 4072 3260 4106 3322
rect 4428 3260 4462 3322
rect 3716 3226 3812 3260
rect 4010 3226 4168 3260
rect 4366 3226 4462 3260
rect -768 2827 -708 2861
rect 3978 2827 4038 2861
rect -768 2801 -734 2827
rect 4004 2801 4038 2827
rect -768 562 -734 588
rect 4004 562 4038 588
rect -768 528 -708 562
rect 3978 528 4038 562
<< psubdiffcont >>
rect 1013 6466 2269 6500
rect 917 5618 951 6404
rect 2331 5618 2365 6404
rect 1013 5522 2269 5556
rect 3292 5536 4432 5570
rect 3196 5336 3230 5474
rect 632 5279 2614 5313
rect 572 3135 606 5253
rect 2640 3135 2674 5253
rect 4494 5336 4528 5474
rect 3292 5240 4432 5274
rect 3808 4766 4407 4800
rect 3748 4300 3782 4740
rect 4433 4300 4467 4740
rect 3808 4240 4407 4274
rect 632 3075 2614 3109
<< nsubdiffcont >>
rect 3812 4078 4010 4112
rect 4168 4078 4366 4112
rect 3716 3322 3750 4016
rect 4072 3322 4106 4016
rect 4428 3322 4462 4016
rect 3812 3226 4010 3260
rect 4168 3226 4366 3260
rect -708 2827 3978 2861
rect -768 588 -734 2801
rect 4004 588 4038 2801
rect -708 528 3978 562
<< poly >>
rect 1003 6324 1091 6340
rect 1003 6056 1019 6324
rect 1053 6056 1091 6324
rect 1003 6040 1091 6056
rect 2191 6324 2279 6340
rect 2191 6056 2229 6324
rect 2263 6056 2279 6324
rect 2191 6040 2279 6056
rect 1003 5966 1091 5982
rect 1003 5698 1019 5966
rect 1053 5698 1091 5966
rect 1003 5682 1091 5698
rect 2191 5966 2279 5982
rect 2191 5698 2229 5966
rect 2263 5698 2279 5966
rect 2191 5682 2279 5698
rect 728 5170 1128 5186
rect 728 5136 744 5170
rect 1112 5136 1128 5170
rect 728 5098 1128 5136
rect 1186 5170 1586 5186
rect 1186 5136 1202 5170
rect 1570 5136 1586 5170
rect 1186 5098 1586 5136
rect 1644 5170 2044 5186
rect 1644 5136 1660 5170
rect 2028 5136 2044 5170
rect 1644 5098 2044 5136
rect 2102 5170 2502 5186
rect 2102 5136 2118 5170
rect 2486 5136 2502 5170
rect 2102 5098 2502 5136
rect 728 4460 1128 4498
rect 728 4426 744 4460
rect 1112 4426 1128 4460
rect 728 4410 1128 4426
rect 1186 4460 1586 4498
rect 1186 4426 1202 4460
rect 1570 4426 1586 4460
rect 1186 4410 1586 4426
rect 1644 4460 2044 4498
rect 1644 4426 1660 4460
rect 2028 4426 2044 4460
rect 1644 4410 2044 4426
rect 2102 4460 2502 4498
rect 2102 4426 2118 4460
rect 2486 4426 2502 4460
rect 2102 4410 2502 4426
rect 728 3963 1128 3979
rect 728 3929 744 3963
rect 1112 3929 1128 3963
rect 728 3891 1128 3929
rect 1186 3963 1586 3979
rect 1186 3929 1202 3963
rect 1570 3929 1586 3963
rect 1186 3891 1586 3929
rect 1644 3963 2044 3979
rect 1644 3929 1660 3963
rect 2028 3929 2044 3963
rect 1644 3891 2044 3929
rect 2102 3963 2502 3979
rect 2102 3929 2118 3963
rect 2486 3929 2502 3963
rect 2102 3891 2502 3929
rect 728 3253 1128 3291
rect 728 3219 744 3253
rect 1112 3219 1128 3253
rect 728 3203 1128 3219
rect 1186 3253 1586 3291
rect 1186 3219 1202 3253
rect 1570 3219 1586 3253
rect 1186 3203 1586 3219
rect 1644 3253 2044 3291
rect 1644 3219 1660 3253
rect 2028 3219 2044 3253
rect 1644 3203 2044 3219
rect 2102 3253 2502 3291
rect 2102 3219 2118 3253
rect 2486 3219 2502 3253
rect 2102 3203 2502 3219
rect 3898 4686 3964 4702
rect 3898 4652 3914 4686
rect 3948 4652 3964 4686
rect 3898 4636 3964 4652
rect 4254 4686 4320 4702
rect 4254 4652 4270 4686
rect 4304 4652 4320 4686
rect 4254 4636 4320 4652
rect 3916 4614 3946 4636
rect 4272 4614 4302 4636
rect 3916 4392 3946 4414
rect 4272 4392 4302 4414
rect 3898 4376 3964 4392
rect 3898 4342 3914 4376
rect 3948 4342 3964 4376
rect 3898 4326 3964 4342
rect 4254 4376 4320 4392
rect 4254 4342 4270 4376
rect 4304 4342 4320 4376
rect 4254 4326 4320 4342
rect 3876 4010 3946 4026
rect 3876 3976 3892 4010
rect 3930 3976 3946 4010
rect 3876 3929 3946 3976
rect 3876 3362 3946 3409
rect 3876 3328 3892 3362
rect 3930 3328 3946 3362
rect 3876 3312 3946 3328
rect 4232 4010 4302 4026
rect 4232 3976 4248 4010
rect 4286 3976 4302 4010
rect 4232 3929 4302 3976
rect 4232 3362 4302 3409
rect 4232 3328 4248 3362
rect 4286 3328 4302 3362
rect 4232 3312 4302 3328
rect -457 2587 543 2603
rect -457 2553 -441 2587
rect 527 2553 543 2587
rect -457 2506 543 2553
rect 601 2587 1601 2603
rect 601 2553 617 2587
rect 1585 2553 1601 2587
rect 601 2506 1601 2553
rect 1659 2587 2659 2603
rect 1659 2553 1675 2587
rect 2643 2553 2659 2587
rect 1659 2506 2659 2553
rect 2717 2587 3717 2603
rect 2717 2553 2733 2587
rect 3701 2553 3717 2587
rect 2717 2506 3717 2553
rect -457 1959 543 2006
rect -457 1925 -441 1959
rect 527 1925 543 1959
rect -457 1909 543 1925
rect 601 1959 1601 2006
rect 601 1925 617 1959
rect 1585 1925 1601 1959
rect 601 1909 1601 1925
rect 1659 1959 2659 2006
rect 1659 1925 1675 1959
rect 2643 1925 2659 1959
rect 1659 1909 2659 1925
rect 2717 1959 3717 2006
rect 2717 1925 2733 1959
rect 3701 1925 3717 1959
rect 2717 1909 3717 1925
rect -457 1425 543 1441
rect -457 1391 -441 1425
rect 527 1391 543 1425
rect -457 1344 543 1391
rect 601 1425 1601 1441
rect 601 1391 617 1425
rect 1585 1391 1601 1425
rect 601 1344 1601 1391
rect 1659 1425 2659 1441
rect 1659 1391 1675 1425
rect 2643 1391 2659 1425
rect 1659 1344 2659 1391
rect 2717 1425 3717 1441
rect 2717 1391 2733 1425
rect 3701 1391 3717 1425
rect 2717 1344 3717 1391
rect -457 797 543 844
rect -457 763 -441 797
rect 527 763 543 797
rect -457 747 543 763
rect 601 797 1601 844
rect 601 763 617 797
rect 1585 763 1601 797
rect 601 747 1601 763
rect 1659 797 2659 844
rect 1659 763 1675 797
rect 2643 763 2659 797
rect 1659 747 2659 763
rect 2717 797 3717 844
rect 2717 763 2733 797
rect 3701 763 3717 797
rect 2717 747 3717 763
<< polycont >>
rect 1019 6056 1053 6324
rect 2229 6056 2263 6324
rect 1019 5698 1053 5966
rect 2229 5698 2263 5966
rect 744 5136 1112 5170
rect 1202 5136 1570 5170
rect 1660 5136 2028 5170
rect 2118 5136 2486 5170
rect 744 4426 1112 4460
rect 1202 4426 1570 4460
rect 1660 4426 2028 4460
rect 2118 4426 2486 4460
rect 744 3929 1112 3963
rect 1202 3929 1570 3963
rect 1660 3929 2028 3963
rect 2118 3929 2486 3963
rect 744 3219 1112 3253
rect 1202 3219 1570 3253
rect 1660 3219 2028 3253
rect 2118 3219 2486 3253
rect 3914 4652 3948 4686
rect 4270 4652 4304 4686
rect 3914 4342 3948 4376
rect 4270 4342 4304 4376
rect 3892 3976 3930 4010
rect 3892 3328 3930 3362
rect 4248 3976 4286 4010
rect 4248 3328 4286 3362
rect -441 2553 527 2587
rect 617 2553 1585 2587
rect 1675 2553 2643 2587
rect 2733 2553 3701 2587
rect -441 1925 527 1959
rect 617 1925 1585 1959
rect 1675 1925 2643 1959
rect 2733 1925 3701 1959
rect -441 1391 527 1425
rect 617 1391 1585 1425
rect 1675 1391 2643 1425
rect 2733 1391 3701 1425
rect -441 763 527 797
rect 617 763 1585 797
rect 1675 763 2643 797
rect 2733 763 3701 797
<< xpolycontact >>
rect 3326 5370 3758 5440
rect 3966 5370 4398 5440
<< xpolyres >>
rect 3758 5370 3966 5440
<< locali >>
rect 494 6770 2647 6821
rect 494 6761 2392 6770
rect 494 5571 503 6761
rect 730 6759 2392 6761
rect 491 5334 503 5571
rect 841 6500 2392 6520
rect 841 6466 1013 6500
rect 2269 6466 2392 6500
rect 841 6441 2392 6466
rect 841 6404 977 6441
rect 841 5618 917 6404
rect 951 5618 977 6404
rect 2331 6404 2392 6441
rect 1087 6352 1103 6386
rect 2179 6352 2195 6386
rect 1019 6324 1053 6340
rect 1019 6040 1053 6056
rect 2229 6324 2263 6340
rect 2229 6040 2263 6056
rect 1087 5994 1103 6028
rect 2179 5994 2195 6028
rect 1019 5966 1053 5982
rect 1019 5682 1053 5698
rect 2229 5966 2263 5982
rect 2229 5682 2263 5698
rect 1087 5636 1103 5670
rect 2179 5636 2195 5670
rect 841 5571 977 5618
rect 2365 5618 2392 6404
rect 2331 5571 2392 5618
rect 841 5556 2392 5571
rect 841 5522 1013 5556
rect 2269 5522 2392 5556
rect 841 5504 2392 5522
rect 2603 5571 2647 6770
rect 2720 5571 4559 5572
rect 2603 5570 4559 5571
rect 2603 5536 3292 5570
rect 4432 5536 4559 5570
rect 2603 5508 4559 5536
rect 2603 5504 3230 5508
rect 3168 5474 3230 5504
rect 3168 5336 3196 5474
rect 4488 5474 4559 5508
rect 491 5233 548 5334
rect 622 5313 2630 5334
rect 622 5279 632 5313
rect 2614 5279 2630 5313
rect 537 4703 548 5233
rect 622 5233 2630 5279
rect 622 4703 630 5233
rect 728 5136 744 5170
rect 1112 5136 1128 5170
rect 1186 5136 1202 5170
rect 1570 5136 1586 5170
rect 1644 5136 1660 5170
rect 2028 5136 2044 5170
rect 2102 5136 2118 5170
rect 2486 5136 2502 5170
rect 537 3667 572 4703
rect 606 3667 630 4703
rect 682 5086 716 5102
rect 682 4494 716 4510
rect 1140 5086 1174 5102
rect 1140 4494 1174 4510
rect 1598 5086 1632 5102
rect 1598 4494 1632 4510
rect 2056 5086 2090 5102
rect 2056 4494 2090 4510
rect 2514 5086 2548 5102
rect 2514 4494 2548 4510
rect 728 4426 744 4460
rect 1112 4426 1128 4460
rect 1186 4426 1202 4460
rect 1570 4426 1586 4460
rect 1644 4426 1660 4460
rect 2028 4426 2044 4460
rect 2102 4426 2118 4460
rect 2486 4426 2502 4460
rect 728 3929 744 3963
rect 1112 3929 1128 3963
rect 1186 3929 1202 3963
rect 1570 3929 1586 3963
rect 1644 3929 1660 3963
rect 2028 3929 2044 3963
rect 2102 3929 2118 3963
rect 2486 3929 2502 3963
rect 537 3151 557 3667
rect 530 3026 557 3151
rect 615 3151 630 3667
rect 682 3879 716 3895
rect 682 3287 716 3303
rect 1140 3879 1174 3895
rect 1140 3287 1174 3303
rect 1598 3879 1632 3895
rect 1598 3287 1632 3303
rect 2056 3879 2090 3895
rect 2056 3287 2090 3303
rect 2514 3879 2548 3895
rect 2514 3287 2548 3303
rect 728 3219 744 3253
rect 1112 3219 1128 3253
rect 1186 3219 1202 3253
rect 1570 3219 1586 3253
rect 1644 3219 1660 3253
rect 2028 3219 2044 3253
rect 2102 3219 2118 3253
rect 2486 3219 2502 3253
rect 2617 3151 2630 5233
rect 615 3129 2630 3151
rect 2706 5232 3048 5334
rect 2706 3123 2739 5232
rect 3025 4886 3048 5232
rect 3168 5296 3230 5336
rect 4488 5336 4494 5474
rect 4528 5336 4559 5474
rect 4488 5296 4559 5336
rect 3168 5274 4559 5296
rect 3168 5240 3292 5274
rect 4432 5240 4559 5274
rect 3168 5158 4559 5240
rect 4426 4886 4559 5158
rect 3025 4800 4559 4886
rect 3025 4766 3808 4800
rect 4407 4766 4559 4800
rect 3025 4749 4559 4766
rect 3025 4740 3800 4749
rect 3025 4300 3748 4740
rect 3782 4300 3800 4740
rect 4413 4740 4559 4749
rect 3898 4652 3914 4686
rect 3948 4652 3964 4686
rect 4254 4652 4270 4686
rect 4304 4652 4320 4686
rect 3870 4602 3904 4618
rect 3870 4410 3904 4426
rect 3958 4602 3992 4618
rect 3958 4410 3992 4426
rect 4226 4602 4260 4618
rect 4226 4410 4260 4426
rect 4314 4602 4348 4618
rect 4314 4410 4348 4426
rect 3898 4342 3914 4376
rect 3948 4342 3964 4376
rect 4254 4342 4270 4376
rect 4304 4342 4320 4376
rect 3025 4298 3800 4300
rect 4413 4300 4433 4740
rect 4467 4300 4559 4740
rect 4413 4298 4559 4300
rect 3025 4274 4559 4298
rect 3025 4240 3808 4274
rect 4407 4240 4559 4274
rect 3025 4220 4559 4240
rect 3623 4112 3761 4135
rect 4424 4112 4507 4121
rect 3623 4078 3812 4112
rect 4010 4078 4168 4112
rect 4366 4078 4507 4112
rect 3623 4052 3761 4078
rect 2706 3026 2731 3123
rect 530 3001 2731 3026
rect 3623 2920 3644 4052
rect 3748 4016 3761 4052
rect 3750 3322 3761 4016
rect 4072 4016 4106 4078
rect 3876 3976 3892 4010
rect 3930 3976 3946 4010
rect 3830 3917 3864 3933
rect 3830 3405 3864 3421
rect 3958 3917 3992 3933
rect 3958 3405 3992 3421
rect 3876 3328 3892 3362
rect 3930 3328 3946 3362
rect -808 2914 3644 2920
rect -822 2893 3644 2914
rect 3748 3279 3761 3322
rect 4424 4016 4507 4078
rect 4232 3976 4248 4010
rect 4286 3976 4302 4010
rect 4186 3917 4220 3933
rect 4186 3405 4220 3421
rect 4314 3917 4348 3933
rect 4314 3405 4348 3421
rect 4232 3328 4248 3362
rect 4286 3328 4302 3362
rect 4072 3279 4106 3322
rect 4424 3322 4428 4016
rect 4462 3322 4507 4016
rect 4424 3279 4507 3322
rect 3748 3260 4507 3279
rect 3748 3226 3812 3260
rect 4010 3226 4168 3260
rect 4366 3226 4507 3260
rect -822 2886 -766 2893
rect -822 706 -801 2886
rect 3748 2861 4507 3226
rect 3978 2838 4507 2861
rect 3978 2827 4120 2838
rect 3748 2801 4120 2827
rect -1013 594 -801 706
rect -1013 229 -863 594
rect 3748 2796 4004 2801
rect -684 2762 4004 2796
rect -684 706 -642 2762
rect -457 2553 -441 2587
rect 527 2553 543 2587
rect 601 2553 617 2587
rect 1585 2553 1601 2587
rect 1659 2553 1675 2587
rect 2643 2553 2659 2587
rect 2717 2553 2733 2587
rect 3701 2553 3717 2587
rect -503 2494 -469 2510
rect -503 2002 -469 2018
rect 555 2494 589 2510
rect 555 2002 589 2018
rect 1613 2494 1647 2510
rect 1613 2002 1647 2018
rect 2671 2494 2705 2510
rect 2671 2002 2705 2018
rect 3729 2494 3763 2510
rect 3729 2002 3763 2018
rect -457 1925 -441 1959
rect 527 1925 543 1959
rect 601 1925 617 1959
rect 1585 1925 1601 1959
rect 1659 1925 1675 1959
rect 2643 1925 2659 1959
rect 2717 1925 2733 1959
rect 3701 1925 3717 1959
rect -457 1391 -441 1425
rect 527 1391 543 1425
rect 601 1391 617 1425
rect 1585 1391 1601 1425
rect 1659 1391 1675 1425
rect 2643 1391 2659 1425
rect 2717 1391 2733 1425
rect 3701 1391 3717 1425
rect 3962 1407 4004 2762
rect 4038 1407 4120 2801
rect -503 1332 -469 1348
rect -503 840 -469 856
rect 555 1332 589 1348
rect 555 840 589 856
rect 1613 1332 1647 1348
rect 1613 840 1647 856
rect 2671 1332 2705 1348
rect 2671 840 2705 856
rect 3729 1332 3763 1348
rect 3729 840 3763 856
rect -457 763 -441 797
rect 527 763 543 797
rect 601 763 617 797
rect 1585 763 1601 797
rect 1659 763 1675 797
rect 2643 763 2659 797
rect 2717 763 2733 797
rect 3701 763 3717 797
rect 3962 706 3983 1407
rect -684 594 3983 706
rect 3941 593 3983 594
rect 4080 593 4120 1407
rect 4099 560 4120 593
rect -1013 228 3840 229
rect 4099 228 4117 560
rect -1013 -144 4117 228
<< viali >>
rect 503 6759 730 6761
rect 2392 6759 2603 6770
rect 503 6520 2603 6759
rect 503 5504 841 6520
rect 1103 6352 2179 6386
rect 1019 6056 1053 6324
rect 2229 6056 2263 6324
rect 1103 5994 2179 6028
rect 1019 5698 1053 5966
rect 2229 5698 2263 5966
rect 1103 5636 2179 5670
rect 2392 5504 2603 6520
rect 503 5334 3168 5504
rect 3344 5386 3741 5424
rect 3983 5386 4380 5424
rect 548 5253 622 5334
rect 548 4703 572 5253
rect 572 4703 606 5253
rect 606 4703 622 5253
rect 2630 5253 2706 5334
rect 744 5136 1112 5170
rect 1202 5136 1570 5170
rect 1660 5136 2028 5170
rect 2118 5136 2486 5170
rect 682 4510 716 5086
rect 1140 4510 1174 5086
rect 1598 4510 1632 5086
rect 2056 4510 2090 5086
rect 2514 4510 2548 5086
rect 744 4426 1112 4460
rect 1202 4426 1570 4460
rect 1660 4426 2028 4460
rect 2118 4426 2486 4460
rect 744 3929 1112 3963
rect 1202 3929 1570 3963
rect 1660 3929 2028 3963
rect 2118 3929 2486 3963
rect 557 3135 572 3667
rect 572 3135 606 3667
rect 606 3135 615 3667
rect 682 3303 716 3879
rect 1140 3303 1174 3879
rect 1598 3303 1632 3879
rect 2056 3303 2090 3879
rect 2514 3303 2548 3879
rect 744 3219 1112 3253
rect 1202 3219 1570 3253
rect 1660 3219 2028 3253
rect 2118 3219 2486 3253
rect 557 3129 615 3135
rect 2630 3135 2640 5253
rect 2640 3135 2674 5253
rect 2674 3135 2706 5253
rect 2630 3129 2706 3135
rect 557 3109 2706 3129
rect 3048 5158 3168 5334
rect 3048 4886 4426 5158
rect 3914 4652 3948 4686
rect 4270 4652 4304 4686
rect 3870 4426 3904 4602
rect 3958 4426 3992 4602
rect 4226 4426 4260 4602
rect 4314 4426 4348 4602
rect 3914 4342 3948 4376
rect 4270 4342 4304 4376
rect 557 3075 632 3109
rect 632 3075 2614 3109
rect 2614 3075 2706 3109
rect 557 3026 2706 3075
rect 3644 4016 3748 4052
rect 3644 3322 3716 4016
rect 3716 3322 3748 4016
rect 3892 3976 3930 4010
rect 3830 3421 3864 3917
rect 3958 3421 3992 3917
rect 3892 3328 3930 3362
rect 3644 2893 3748 3322
rect 4248 3976 4286 4010
rect 4186 3421 4220 3917
rect 4314 3421 4348 3917
rect 4248 3328 4286 3362
rect -766 2886 3748 2893
rect -801 2861 3748 2886
rect -801 2827 -708 2861
rect -708 2827 3748 2861
rect -801 2801 3748 2827
rect -801 594 -768 2801
rect -863 588 -768 594
rect -768 588 -734 2801
rect -734 2796 3748 2801
rect -734 594 -684 2796
rect -441 2553 527 2587
rect 617 2553 1585 2587
rect 1675 2553 2643 2587
rect 2733 2553 3701 2587
rect -503 2018 -469 2494
rect 555 2018 589 2494
rect 1613 2018 1647 2494
rect 2671 2018 2705 2494
rect 3729 2018 3763 2494
rect -441 1925 527 1959
rect 617 1925 1585 1959
rect 1675 1925 2643 1959
rect 2733 1925 3701 1959
rect -441 1391 527 1425
rect 617 1391 1585 1425
rect 1675 1391 2643 1425
rect 2733 1391 3701 1425
rect -503 856 -469 1332
rect 555 856 589 1332
rect 1613 856 1647 1332
rect 2671 856 2705 1332
rect 3729 856 3763 1332
rect -441 763 527 797
rect 617 763 1585 797
rect 1675 763 2643 797
rect 2733 763 3701 797
rect -734 593 3941 594
rect 3983 593 4004 1407
rect -734 588 4004 593
rect 4004 588 4038 1407
rect 4038 593 4080 1407
rect 4038 588 4099 593
rect -863 562 4099 588
rect -863 528 -708 562
rect -708 528 3978 562
rect 3978 528 4099 562
rect -863 229 4099 528
rect 3840 228 4099 229
<< metal1 >>
rect 497 6765 736 6773
rect 2386 6770 2609 6782
rect 2382 6765 2392 6770
rect 497 6761 2392 6765
rect 493 5334 503 6761
rect 730 6759 2392 6761
rect 841 6514 2392 6520
rect 841 5511 851 6514
rect 1760 6392 1770 6401
rect 1091 6386 1770 6392
rect 2179 6392 2189 6401
rect 1091 6352 1103 6386
rect 1091 6346 1770 6352
rect 1760 6336 1770 6346
rect 2179 6346 2191 6392
rect 2179 6336 2189 6346
rect 1013 6324 1059 6336
rect 1013 6056 1019 6324
rect 1053 6056 1059 6324
rect 1013 5966 1059 6056
rect 2223 6324 2269 6336
rect 2223 6056 2229 6324
rect 2263 6056 2269 6324
rect 1093 6034 1103 6043
rect 1091 5988 1103 6034
rect 1603 6034 1613 6043
rect 1603 6028 2191 6034
rect 2179 5994 2191 6028
rect 1093 5979 1103 5988
rect 1603 5988 2191 5994
rect 1603 5979 1613 5988
rect 1013 5853 1019 5966
rect 1053 5853 1059 5966
rect 2223 5966 2269 6056
rect 998 5713 1008 5853
rect 1064 5713 1074 5853
rect 1013 5698 1019 5713
rect 1053 5698 1059 5713
rect 1013 5686 1059 5698
rect 2223 5698 2229 5966
rect 2263 5698 2269 5966
rect 2223 5686 2269 5698
rect 1760 5676 1770 5685
rect 1091 5670 1770 5676
rect 2179 5676 2189 5685
rect 1091 5636 1103 5670
rect 1091 5630 1770 5636
rect 1760 5620 1770 5630
rect 2179 5630 2191 5676
rect 2179 5620 2189 5630
rect 1846 5510 1856 5511
rect 2382 5510 2392 6514
rect 1846 5504 2392 5510
rect 2603 5510 2613 6770
rect 2973 5510 3174 5516
rect 2603 5504 3174 5510
rect 497 5322 548 5334
rect 538 4703 548 5322
rect 622 5328 2630 5334
rect 622 5322 736 5328
rect 622 4703 632 5322
rect 732 5170 1124 5176
rect 732 5136 744 5170
rect 1112 5136 1124 5170
rect 732 5130 1124 5136
rect 1190 5170 1582 5176
rect 1190 5136 1202 5170
rect 1570 5136 1582 5170
rect 1190 5130 1582 5136
rect 1648 5170 2040 5176
rect 1648 5136 1660 5170
rect 2028 5136 2040 5170
rect 1648 5130 2040 5136
rect 2106 5170 2498 5176
rect 2106 5136 2118 5170
rect 2486 5136 2498 5170
rect 2106 5130 2498 5136
rect 676 5086 722 5098
rect 1134 5086 1180 5098
rect 1592 5086 1638 5098
rect 2050 5086 2096 5098
rect 2508 5086 2554 5098
rect 542 4691 628 4703
rect 676 4658 682 5086
rect 716 4658 722 5086
rect 1121 4926 1131 5086
rect 1183 4926 1193 5086
rect 641 4521 651 4658
rect 745 4521 755 4658
rect 676 4510 682 4521
rect 716 4510 722 4521
rect 676 4498 722 4510
rect 1134 4510 1140 4926
rect 1174 4510 1180 4926
rect 1592 4869 1598 5086
rect 1632 4869 1638 5086
rect 2037 4926 2047 5086
rect 2099 4926 2109 5086
rect 1558 4732 1568 4869
rect 1662 4732 1672 4869
rect 1134 4498 1180 4510
rect 1592 4510 1598 4732
rect 1632 4510 1638 4732
rect 1592 4498 1638 4510
rect 2050 4510 2056 4926
rect 2090 4510 2096 4926
rect 2508 4658 2514 5086
rect 2548 4658 2554 5086
rect 2473 4521 2483 4658
rect 2577 4521 2587 4658
rect 2050 4498 2096 4510
rect 2508 4510 2514 4521
rect 2548 4510 2554 4521
rect 2508 4498 2554 4510
rect 734 4466 744 4469
rect 732 4420 744 4466
rect 944 4466 954 4469
rect 1192 4466 1202 4469
rect 944 4460 1124 4466
rect 1112 4426 1124 4460
rect 734 4417 744 4420
rect 944 4420 1124 4426
rect 1190 4420 1202 4466
rect 1402 4466 1412 4469
rect 1650 4466 1660 4469
rect 1402 4460 1582 4466
rect 1570 4426 1582 4460
rect 944 4417 954 4420
rect 1192 4417 1202 4420
rect 1402 4420 1582 4426
rect 1648 4420 1660 4466
rect 1860 4466 1870 4469
rect 2108 4466 2118 4469
rect 1860 4460 2040 4466
rect 2028 4426 2040 4460
rect 1402 4417 1412 4420
rect 1650 4417 1660 4420
rect 1860 4420 2040 4426
rect 2106 4420 2118 4466
rect 2318 4466 2328 4469
rect 2318 4460 2498 4466
rect 2486 4426 2498 4460
rect 1860 4417 1870 4420
rect 2108 4417 2118 4420
rect 2318 4420 2498 4426
rect 2318 4417 2328 4420
rect -67 4230 744 4330
rect 844 4230 1470 4330
rect 1570 4230 1928 4330
rect 2028 4230 2118 4330
rect 2218 4230 2531 4330
rect -67 4044 1012 4144
rect 1112 4044 1202 4144
rect 1302 4044 1660 4144
rect 1760 4044 2386 4144
rect 2486 4044 2531 4144
rect 902 3969 912 3972
rect 732 3963 912 3969
rect 1112 3969 1122 3972
rect 1360 3969 1370 3972
rect 732 3929 744 3963
rect 732 3923 912 3929
rect 902 3920 912 3923
rect 1112 3923 1124 3969
rect 1190 3963 1370 3969
rect 1570 3969 1580 3972
rect 1818 3969 1828 3972
rect 1190 3929 1202 3963
rect 1190 3923 1370 3929
rect 1112 3920 1122 3923
rect 1360 3920 1370 3923
rect 1570 3923 1582 3969
rect 1648 3963 1828 3969
rect 2028 3969 2038 3972
rect 2276 3969 2286 3972
rect 1648 3929 1660 3963
rect 1648 3923 1828 3929
rect 1570 3920 1580 3923
rect 1818 3920 1828 3923
rect 2028 3923 2040 3969
rect 2106 3963 2286 3969
rect 2486 3969 2496 3972
rect 2106 3929 2118 3963
rect 2106 3923 2286 3929
rect 2028 3920 2038 3923
rect 2276 3920 2286 3923
rect 2486 3923 2498 3969
rect 2486 3920 2496 3923
rect 676 3879 722 3891
rect 676 3869 682 3879
rect 716 3869 722 3879
rect 1134 3879 1180 3891
rect 640 3732 650 3869
rect 744 3732 754 3869
rect 551 3667 621 3679
rect 547 3026 557 3667
rect 615 3135 625 3667
rect 676 3303 682 3732
rect 716 3303 722 3732
rect 1134 3463 1140 3879
rect 1174 3463 1180 3879
rect 1592 3879 1638 3891
rect 1592 3611 1598 3879
rect 1632 3611 1638 3879
rect 2050 3879 2096 3891
rect 1559 3474 1569 3611
rect 1663 3474 1673 3611
rect 1121 3303 1131 3463
rect 1183 3303 1193 3463
rect 1592 3303 1598 3474
rect 1632 3303 1638 3474
rect 2050 3463 2056 3879
rect 2090 3463 2096 3879
rect 2508 3879 2554 3891
rect 2508 3869 2514 3879
rect 2548 3869 2554 3879
rect 2475 3732 2485 3869
rect 2579 3732 2589 3869
rect 2037 3303 2047 3463
rect 2099 3303 2109 3463
rect 2508 3303 2514 3732
rect 2548 3303 2554 3732
rect 676 3291 722 3303
rect 1134 3291 1180 3303
rect 1592 3291 1638 3303
rect 2050 3291 2096 3303
rect 2508 3291 2554 3303
rect 732 3253 1124 3259
rect 732 3219 744 3253
rect 1112 3219 1124 3253
rect 732 3213 1124 3219
rect 1190 3253 1582 3259
rect 1190 3219 1202 3253
rect 1570 3219 1582 3253
rect 1190 3213 1582 3219
rect 1648 3253 2040 3259
rect 1648 3219 1660 3253
rect 2028 3219 2040 3253
rect 1648 3213 2040 3219
rect 2106 3253 2498 3259
rect 2106 3219 2118 3253
rect 2486 3219 2498 3253
rect 2106 3213 2498 3219
rect 2624 3135 2630 5328
rect 615 3129 2630 3135
rect 2706 5328 3048 5334
rect 2706 3026 2712 5328
rect 2973 5322 3048 5328
rect 3042 5164 3048 5322
rect 3036 4886 3048 5164
rect 3168 5164 3174 5504
rect 4168 5430 4178 5431
rect 3332 5380 3344 5430
rect 3546 5424 3753 5430
rect 3741 5386 3753 5424
rect 3334 5378 3344 5380
rect 3546 5380 3753 5386
rect 3971 5424 4178 5430
rect 4380 5430 4390 5431
rect 3971 5386 3983 5424
rect 3971 5380 4178 5386
rect 3546 5378 3556 5380
rect 4168 5379 4178 5380
rect 4380 5380 4392 5430
rect 4380 5379 4390 5380
rect 3168 5158 4438 5164
rect 4426 4886 4438 5158
rect 3036 4880 4438 4886
rect 3902 4686 4316 4692
rect 3902 4652 3914 4686
rect 3948 4652 4270 4686
rect 4304 4652 4316 4686
rect 3902 4646 4316 4652
rect 3864 4602 3910 4614
rect 3952 4602 3998 4614
rect 4220 4602 4266 4614
rect 4308 4602 4354 4614
rect 3851 4531 3861 4602
rect 3913 4531 3923 4602
rect 3864 4426 3870 4531
rect 3904 4426 3910 4531
rect 3864 4414 3910 4426
rect 3952 4426 3958 4602
rect 3992 4426 3998 4602
rect 4207 4531 4217 4602
rect 4269 4531 4279 4602
rect 3952 4414 3998 4426
rect 4220 4426 4226 4531
rect 4260 4426 4266 4531
rect 4308 4497 4314 4602
rect 4348 4497 4354 4602
rect 4295 4426 4305 4497
rect 4357 4426 4367 4497
rect 4220 4414 4266 4426
rect 4308 4414 4354 4426
rect 3958 4382 3992 4414
rect 3902 4376 3949 4382
rect 3902 4342 3914 4376
rect 3948 4342 3949 4376
rect 3902 4336 3949 4342
rect 3939 4303 3949 4336
rect 4001 4376 4316 4382
rect 4001 4342 4270 4376
rect 4304 4342 4316 4376
rect 4001 4336 4316 4342
rect 4001 4303 4011 4336
rect 3638 4052 3754 4064
rect 551 3020 2712 3026
rect 551 3014 621 3020
rect 2624 3014 2712 3020
rect 3634 2899 3644 4052
rect -778 2898 3644 2899
rect -807 2893 3644 2898
rect 3748 2899 3758 4052
rect 3878 4010 3943 4027
rect 3878 3976 3892 4010
rect 3930 3976 3943 4010
rect 3878 3969 3943 3976
rect 4236 4010 4298 4041
rect 4236 3976 4248 4010
rect 4286 3976 4298 4010
rect 4236 3970 4298 3976
rect 3824 3917 3870 3929
rect 3952 3917 3998 3929
rect 4180 3917 4226 3929
rect 4308 3917 4354 3929
rect 3824 3621 3830 3917
rect 3864 3621 3870 3917
rect 3939 3717 3949 3917
rect 4001 3717 4011 3917
rect 3811 3421 3821 3621
rect 3873 3421 3883 3621
rect 3952 3421 3958 3717
rect 3992 3421 3998 3717
rect 4180 3621 4186 3917
rect 4220 3621 4226 3917
rect 4295 3717 4305 3917
rect 4357 3717 4367 3917
rect 4167 3421 4177 3621
rect 4229 3421 4239 3621
rect 4308 3421 4314 3717
rect 4348 3421 4354 3717
rect 3824 3409 3870 3421
rect 3952 3409 3998 3421
rect 4180 3409 4226 3421
rect 4308 3409 4354 3421
rect 3861 3362 3961 3368
rect 3861 3328 3892 3362
rect 3930 3328 3961 3362
rect -807 2886 -766 2893
rect -811 600 -801 2886
rect 3748 2796 3760 2899
rect -875 594 -801 600
rect -684 2790 3760 2796
rect -684 600 -674 2790
rect -509 2587 539 2593
rect -509 2553 -441 2587
rect 527 2553 539 2587
rect -509 2547 539 2553
rect 605 2587 2655 2593
rect 605 2553 617 2587
rect 1585 2553 1675 2587
rect 2643 2553 2655 2587
rect 605 2547 2655 2553
rect 2721 2587 3769 2593
rect 2721 2553 2733 2587
rect 3701 2553 3769 2587
rect 2721 2547 3769 2553
rect -509 2494 -463 2547
rect 549 2494 595 2506
rect 1607 2494 1653 2547
rect 2665 2494 2711 2506
rect 3723 2494 3769 2547
rect -509 2218 -503 2494
rect -469 2218 -463 2494
rect -528 2018 -518 2218
rect -454 2018 -444 2218
rect 536 2194 546 2494
rect 598 2194 608 2494
rect 1588 2294 1598 2494
rect 1662 2294 1672 2494
rect 549 2018 555 2194
rect 589 2018 595 2194
rect -509 1969 -463 2018
rect 549 2006 595 2018
rect 1607 2018 1613 2294
rect 1647 2018 1653 2294
rect 2652 2194 2662 2494
rect 2714 2194 2724 2494
rect 3723 2218 3729 2494
rect 3763 2218 3769 2494
rect -509 1968 -431 1969
rect 1607 1968 1653 2018
rect 2665 2018 2671 2194
rect 2705 2018 2711 2194
rect 3704 2018 3714 2218
rect 3778 2018 3788 2218
rect 2665 2006 2711 2018
rect -509 1916 -441 1968
rect 199 1965 209 1968
rect 607 1965 617 1968
rect 199 1959 539 1965
rect 527 1925 539 1959
rect 199 1919 539 1925
rect 605 1919 617 1965
rect 1257 1965 1267 1968
rect 1607 1965 1675 1968
rect 1257 1959 1675 1965
rect 2315 1965 2325 1968
rect 2723 1965 2733 1968
rect 2315 1959 2655 1965
rect 1585 1925 1675 1959
rect 2643 1925 2655 1959
rect 199 1916 209 1919
rect 607 1916 617 1919
rect 1257 1919 1675 1925
rect 1257 1916 1267 1919
rect 1665 1916 1675 1919
rect 2315 1919 2655 1925
rect 2721 1919 2733 1965
rect 3373 1965 3383 1968
rect 3723 1965 3769 2018
rect 3373 1959 3769 1965
rect 3701 1925 3769 1959
rect 2315 1916 2325 1919
rect 2723 1916 2733 1919
rect 3373 1919 3769 1925
rect 3373 1916 3383 1919
rect -509 1915 -463 1916
rect 3861 1812 3961 3328
rect -457 1712 -441 1812
rect -341 1712 1485 1812
rect 1585 1712 2543 1812
rect 2643 1712 2733 1812
rect 2833 1712 3961 1812
rect 4216 3362 4316 3368
rect 4216 3328 4248 3362
rect 4286 3328 4316 3362
rect 4216 1630 4316 3328
rect -460 1530 427 1630
rect 527 1530 617 1630
rect 717 1530 1675 1630
rect 1775 1530 3601 1630
rect 3701 1530 4316 1630
rect -123 1431 -113 1434
rect -509 1425 -113 1431
rect 527 1431 537 1434
rect 935 1431 945 1434
rect -509 1391 -441 1425
rect -509 1385 -113 1391
rect -509 1332 -463 1385
rect -123 1382 -113 1385
rect 527 1385 539 1431
rect 605 1425 945 1431
rect 1585 1431 1668 1434
rect 1993 1431 2003 1433
rect 1585 1425 2003 1431
rect 2643 1431 2653 1433
rect 3051 1431 3061 1434
rect 605 1391 617 1425
rect 1585 1391 1675 1425
rect 605 1385 945 1391
rect 527 1382 537 1385
rect 935 1382 945 1385
rect 1585 1385 2003 1391
rect 1585 1382 1668 1385
rect 549 1332 595 1344
rect -528 1132 -518 1332
rect -454 1132 -444 1332
rect 549 1156 555 1332
rect 589 1156 595 1332
rect 1607 1332 1653 1382
rect 1993 1381 2003 1385
rect 2643 1385 2655 1431
rect 2721 1425 3061 1431
rect 3701 1431 3711 1434
rect 2721 1391 2733 1425
rect 2721 1385 3061 1391
rect 2643 1381 2653 1385
rect 3051 1382 3061 1385
rect 3701 1385 3713 1431
rect 3977 1407 4086 1419
rect 3701 1382 3711 1385
rect -509 856 -503 1132
rect -469 856 -463 1132
rect 536 856 546 1156
rect 598 856 608 1156
rect 1607 1056 1613 1332
rect 1647 1056 1653 1332
rect 2665 1332 2711 1344
rect 3723 1332 3769 1344
rect 2665 1156 2671 1332
rect 2705 1156 2711 1332
rect 1588 856 1598 1056
rect 1662 856 1672 1056
rect 2652 856 2662 1156
rect 2714 856 2724 1156
rect 3704 1132 3714 1332
rect 3778 1132 3788 1332
rect 3723 856 3729 1132
rect 3763 856 3769 1132
rect -509 803 -463 856
rect 549 844 595 856
rect 1607 803 1653 856
rect 2665 844 2711 856
rect 3723 803 3769 856
rect -509 797 539 803
rect -509 763 -441 797
rect 527 763 539 797
rect -509 757 539 763
rect 605 797 2655 803
rect 605 763 617 797
rect 1585 763 1675 797
rect 2643 763 2655 797
rect 605 757 2655 763
rect 2721 797 3769 803
rect 2721 763 2733 797
rect 3701 763 3769 797
rect 2721 757 3769 763
rect 3973 605 3983 1407
rect 3834 600 3983 605
rect -684 594 3983 600
rect -875 229 -863 594
rect 3941 593 3983 594
rect 4080 605 4090 1407
rect 4080 593 4105 605
rect -875 228 3840 229
rect 4099 228 4109 593
rect -875 223 4105 228
rect 3834 216 4105 223
<< via1 >>
rect 503 6759 730 6761
rect 2392 6759 2603 6770
rect 503 6520 2603 6759
rect 503 5504 841 6520
rect 1770 6386 2179 6401
rect 1770 6352 2179 6386
rect 1770 6336 2179 6352
rect 1103 6028 1603 6043
rect 1103 5994 1603 6028
rect 1103 5979 1603 5994
rect 1008 5713 1019 5853
rect 1019 5713 1053 5853
rect 1053 5713 1064 5853
rect 1770 5670 2179 5685
rect 1770 5636 2179 5670
rect 1770 5620 2179 5636
rect 841 5504 1846 5511
rect 503 5341 1846 5504
rect 2392 5469 2603 6520
rect 503 5334 730 5341
rect 548 4703 622 5334
rect 1131 4926 1140 5086
rect 1140 4926 1174 5086
rect 1174 4926 1183 5086
rect 651 4521 682 4658
rect 682 4521 716 4658
rect 716 4521 745 4658
rect 2047 4926 2056 5086
rect 2056 4926 2090 5086
rect 2090 4926 2099 5086
rect 1568 4732 1598 4869
rect 1598 4732 1632 4869
rect 1632 4732 1662 4869
rect 2483 4521 2514 4658
rect 2514 4521 2548 4658
rect 2548 4521 2577 4658
rect 744 4460 944 4469
rect 744 4426 944 4460
rect 744 4417 944 4426
rect 1202 4460 1402 4469
rect 1202 4426 1402 4460
rect 1202 4417 1402 4426
rect 1660 4460 1860 4469
rect 1660 4426 1860 4460
rect 1660 4417 1860 4426
rect 2118 4460 2318 4469
rect 2118 4426 2318 4460
rect 2118 4417 2318 4426
rect 744 4230 844 4330
rect 1470 4230 1570 4330
rect 1928 4230 2028 4330
rect 2118 4230 2218 4330
rect 1012 4044 1112 4144
rect 1202 4044 1302 4144
rect 1660 4044 1760 4144
rect 2386 4044 2486 4144
rect 912 3963 1112 3972
rect 912 3929 1112 3963
rect 912 3920 1112 3929
rect 1370 3963 1570 3972
rect 1370 3929 1570 3963
rect 1370 3920 1570 3929
rect 1828 3963 2028 3972
rect 1828 3929 2028 3963
rect 1828 3920 2028 3929
rect 2286 3963 2486 3972
rect 2286 3929 2486 3963
rect 2286 3920 2486 3929
rect 650 3732 682 3869
rect 682 3732 716 3869
rect 716 3732 744 3869
rect 557 3129 615 3667
rect 1569 3474 1598 3611
rect 1598 3474 1632 3611
rect 1632 3474 1663 3611
rect 1131 3303 1140 3463
rect 1140 3303 1174 3463
rect 1174 3303 1183 3463
rect 2485 3732 2514 3869
rect 2514 3732 2548 3869
rect 2548 3732 2579 3869
rect 2047 3303 2056 3463
rect 2056 3303 2090 3463
rect 2090 3303 2099 3463
rect 557 3026 2685 3129
rect 3344 5424 3546 5430
rect 3344 5386 3546 5424
rect 3344 5378 3546 5386
rect 4178 5424 4380 5431
rect 4178 5386 4380 5424
rect 4178 5379 4380 5386
rect 3048 4886 4426 5158
rect 3861 4531 3870 4602
rect 3870 4531 3904 4602
rect 3904 4531 3913 4602
rect 4217 4531 4226 4602
rect 4226 4531 4260 4602
rect 4260 4531 4269 4602
rect 4305 4426 4314 4497
rect 4314 4426 4348 4497
rect 4348 4426 4357 4497
rect 3949 4303 4001 4382
rect 3644 2893 3748 4052
rect 3949 3717 3958 3917
rect 3958 3717 3992 3917
rect 3992 3717 4001 3917
rect 3821 3421 3830 3621
rect 3830 3421 3864 3621
rect 3864 3421 3873 3621
rect 4305 3717 4314 3917
rect 4314 3717 4348 3917
rect 4348 3717 4357 3917
rect 4177 3421 4186 3621
rect 4186 3421 4220 3621
rect 4220 3421 4229 3621
rect -766 2886 3748 2893
rect -801 2796 3748 2886
rect -801 594 -684 2796
rect -518 2018 -503 2218
rect -503 2018 -469 2218
rect -469 2018 -454 2218
rect 546 2194 555 2494
rect 555 2194 589 2494
rect 589 2194 598 2494
rect 1598 2294 1613 2494
rect 1613 2294 1647 2494
rect 1647 2294 1662 2494
rect 2662 2194 2671 2494
rect 2671 2194 2705 2494
rect 2705 2194 2714 2494
rect 3714 2018 3729 2218
rect 3729 2018 3763 2218
rect 3763 2018 3778 2218
rect -441 1959 199 1968
rect -441 1925 199 1959
rect -441 1916 199 1925
rect 617 1959 1257 1968
rect 1675 1959 2315 1968
rect 617 1925 1257 1959
rect 1675 1925 2315 1959
rect 617 1916 1257 1925
rect 1675 1916 2315 1925
rect 2733 1959 3373 1968
rect 2733 1925 3373 1959
rect 2733 1916 3373 1925
rect -441 1712 -341 1812
rect 1485 1712 1585 1812
rect 2543 1712 2643 1812
rect 2733 1712 2833 1812
rect 427 1530 527 1630
rect 617 1530 717 1630
rect 1675 1530 1775 1630
rect 3601 1530 3701 1630
rect -113 1425 527 1434
rect -113 1391 527 1425
rect -113 1382 527 1391
rect 945 1425 1585 1434
rect 2003 1425 2643 1433
rect 945 1391 1585 1425
rect 2003 1391 2643 1425
rect 945 1382 1585 1391
rect -518 1132 -503 1332
rect -503 1132 -469 1332
rect -469 1132 -454 1332
rect 2003 1381 2643 1391
rect 3061 1425 3701 1434
rect 3061 1391 3701 1425
rect 3061 1382 3701 1391
rect 546 856 555 1156
rect 555 856 589 1156
rect 589 856 598 1156
rect 1598 856 1613 1056
rect 1613 856 1647 1056
rect 1647 856 1662 1056
rect 2662 856 2671 1156
rect 2671 856 2705 1156
rect 2705 856 2714 1156
rect 3714 1132 3729 1332
rect 3729 1132 3763 1332
rect 3763 1132 3778 1332
rect -863 593 3941 594
rect 3983 593 4080 1407
rect -863 229 4099 593
rect 3840 228 4099 229
<< metal2 >>
rect 461 6771 621 6772
rect 461 6769 730 6771
rect 2392 6770 2603 6780
rect 461 6761 2392 6769
rect 461 6487 503 6761
rect 730 6759 2392 6761
rect 841 6510 2392 6520
rect 1770 6401 2179 6411
rect 1770 6326 2179 6336
rect 841 6043 1603 6053
rect 841 5979 1103 6043
rect 841 5969 1603 5979
rect 1008 5853 1064 5863
rect 1008 5703 1064 5713
rect 2056 5695 2178 6326
rect 1770 5685 2179 5695
rect 1770 5610 2179 5620
rect 841 5511 1846 5521
rect 730 5334 1846 5341
rect 503 5324 548 5334
rect 622 5331 1846 5334
rect 622 5324 730 5331
rect 2056 5096 2178 5610
rect 2392 5459 2603 5469
rect 3138 5430 3279 5440
rect 3344 5430 3546 5440
rect 3279 5378 3344 5430
rect 3279 5368 3546 5378
rect 4178 5431 4660 5441
rect 4380 5379 4660 5431
rect 4178 5369 4660 5379
rect 3138 5358 3279 5368
rect 1131 5093 1183 5096
rect 2047 5093 2178 5096
rect 3048 5158 4426 5168
rect 1131 5086 2979 5093
rect 1183 4993 2047 5086
rect 1131 4916 1183 4926
rect 2099 4993 2979 5086
rect 2047 4916 2099 4926
rect 1568 4869 1662 4879
rect 1568 4722 1662 4732
rect 548 4693 622 4703
rect 651 4658 745 4668
rect 651 4511 745 4521
rect 2483 4658 2577 4668
rect 2483 4511 2577 4521
rect 744 4469 944 4479
rect 744 4407 944 4417
rect 1202 4469 1402 4479
rect 1202 4407 1402 4417
rect 1660 4469 1860 4479
rect 1660 4407 1860 4417
rect 2118 4469 2318 4479
rect 2118 4407 2318 4417
rect 744 4330 844 4407
rect 744 4220 844 4230
rect 1012 4144 1112 4154
rect 1012 3982 1112 4044
rect 1202 4144 1302 4407
rect 1202 4034 1302 4044
rect 1470 4330 1570 4340
rect 1470 3982 1570 4230
rect 1660 4144 1760 4407
rect 1660 4034 1760 4044
rect 1928 4330 2028 4340
rect 1928 3982 2028 4230
rect 2118 4330 2218 4407
rect 2118 4220 2218 4230
rect 2386 4144 2486 4154
rect 2386 3982 2486 4044
rect 912 3972 1112 3982
rect 912 3910 1112 3920
rect 1370 3972 1570 3982
rect 1370 3910 1570 3920
rect 1828 3972 2028 3982
rect 1828 3910 2028 3920
rect 2286 3972 2486 3982
rect 2286 3910 2486 3920
rect 650 3869 744 3879
rect 650 3722 744 3732
rect 2485 3869 2579 3879
rect 2485 3722 2579 3732
rect 557 3667 615 3677
rect 1569 3611 1663 3621
rect 1131 3463 1183 3473
rect 1569 3464 1663 3474
rect 2047 3463 2099 3473
rect 1183 3303 2047 3394
rect 2879 3394 2979 4993
rect 3048 4876 4426 4886
rect 3861 4602 3913 4876
rect 3861 4521 3913 4531
rect 4217 4602 4269 4876
rect 4217 4521 4269 4531
rect 4305 4497 4357 4507
rect 3949 4382 4001 4392
rect 2099 3303 2979 3394
rect 1131 3294 2979 3303
rect 3644 4052 3748 4062
rect 1131 3293 1183 3294
rect 2047 3293 2099 3294
rect 615 3129 2685 3139
rect 557 3016 2685 3026
rect -766 2896 3644 2903
rect -801 2893 3644 2896
rect 3949 3917 4001 4303
rect 3949 3707 4001 3717
rect 4305 4253 4357 4426
rect 4588 4253 4660 5369
rect 4305 4181 4779 4253
rect 4305 3917 4357 4181
rect 4305 3707 4357 3717
rect 3821 3621 3873 3631
rect 3748 3421 3821 3553
rect 4177 3621 4229 3631
rect 3873 3421 4177 3553
rect 3748 3411 4229 3421
rect -801 2886 -766 2893
rect -863 594 -801 604
rect -684 2786 3748 2796
rect 546 2494 598 2786
rect -518 2218 -454 2228
rect 1598 2494 1662 2504
rect 1598 2284 1662 2294
rect 2662 2494 2714 2786
rect 546 2184 598 2194
rect 2662 2184 2714 2194
rect 3714 2218 3778 2228
rect -518 2008 -454 2018
rect 3714 2008 3778 2018
rect -441 1968 199 1978
rect -441 1906 199 1916
rect 617 1968 1257 1978
rect 617 1906 1257 1916
rect 1675 1968 2315 1978
rect 1675 1906 2315 1916
rect 2733 1968 3373 1978
rect 2733 1906 3373 1916
rect -441 1812 -341 1906
rect -441 1702 -341 1712
rect 427 1630 527 1640
rect 427 1444 527 1530
rect 617 1630 717 1906
rect 617 1520 717 1530
rect 1485 1812 1585 1822
rect 1485 1444 1585 1712
rect 1675 1630 1775 1906
rect 1675 1520 1775 1530
rect 2543 1812 2643 1822
rect -113 1434 527 1444
rect -113 1372 527 1382
rect 945 1434 1585 1444
rect 2543 1443 2643 1712
rect 2733 1812 2833 1906
rect 2733 1702 2833 1712
rect 3601 1630 3701 1640
rect 3601 1444 3701 1530
rect 945 1372 1585 1382
rect 2003 1433 2643 1443
rect 2003 1371 2643 1381
rect 3061 1434 3701 1444
rect 3061 1372 3701 1382
rect 3983 1407 4080 1417
rect -518 1332 -454 1342
rect 3714 1332 3778 1342
rect -518 1122 -454 1132
rect 546 1156 598 1166
rect 2662 1156 2714 1166
rect 546 604 598 856
rect 1598 1056 1662 1066
rect 1598 846 1662 856
rect 3714 1122 3778 1132
rect 2662 604 2714 856
rect -684 603 3941 604
rect -684 594 3983 603
rect 3941 593 3983 594
rect 4080 602 4099 603
rect 4080 593 4217 602
rect -863 228 3840 229
rect 4099 228 4217 593
rect -863 219 4217 228
rect 3840 218 4217 219
rect 4079 217 4217 218
<< via2 >>
rect 1008 5713 1064 5853
rect 3138 5368 3279 5430
rect 1568 4732 1662 4869
rect 651 4521 745 4658
rect 2483 4521 2577 4658
rect 650 3732 744 3869
rect 2485 3732 2579 3869
rect 1569 3474 1663 3611
rect -518 2018 -454 2218
rect 1598 2294 1662 2494
rect 3714 2018 3778 2218
rect -518 1132 -454 1332
rect 1598 856 1662 1056
rect 3714 1132 3778 1332
<< metal3 >>
rect 2840 9406 6612 9434
rect 2840 7034 6528 9406
rect 2618 6927 6528 7034
rect 2840 5982 6528 6927
rect 6592 5982 6612 9406
rect 2840 5954 6612 5982
rect 998 5853 1074 5858
rect 998 5768 1008 5853
rect 220 5713 1008 5768
rect 1064 5713 1074 5853
rect 220 5708 1074 5713
rect 220 4563 280 5708
rect 3128 5433 3289 5435
rect 3128 5365 3138 5433
rect 3279 5365 3289 5433
rect 3128 5363 3289 5365
rect 1558 4869 2905 4874
rect 1558 4732 1568 4869
rect 1662 4732 2905 4869
rect 1558 4727 1672 4732
rect -67 4503 280 4563
rect 641 4658 755 4663
rect 641 4521 651 4658
rect 745 4521 755 4658
rect 641 4516 755 4521
rect 2473 4658 2587 4663
rect 2473 4521 2483 4658
rect 2577 4521 2587 4658
rect 2473 4516 2587 4521
rect 2758 3874 2905 4732
rect 640 3869 2905 3874
rect 640 3732 650 3869
rect 744 3732 2485 3869
rect 2579 3732 2905 3869
rect 640 3727 2905 3732
rect 1559 3611 1673 3616
rect 1559 3474 1569 3611
rect 1663 3474 1673 3611
rect 1559 3469 1673 3474
rect 2758 2499 2905 3727
rect 1588 2494 4228 2499
rect 1588 2294 1598 2494
rect 1662 2399 4228 2494
rect 1662 2294 1672 2399
rect 1588 2289 1672 2294
rect -528 2218 -444 2223
rect -528 2018 -518 2218
rect -454 2018 -444 2218
rect -528 2013 -444 2018
rect 3704 2218 3788 2223
rect 3704 2018 3714 2218
rect 3778 2018 3788 2218
rect 3704 2013 3788 2018
rect 4128 1337 4228 2399
rect -528 1332 4228 1337
rect -528 1132 -518 1332
rect -454 1237 3714 1332
rect -454 1132 -444 1237
rect -528 1127 -444 1132
rect 3704 1132 3714 1237
rect 3778 1237 4228 1332
rect 3778 1132 3788 1237
rect 3704 1127 3788 1132
rect 1588 1056 1672 1061
rect 1588 856 1598 1056
rect 1662 856 1672 1056
rect 1588 851 1672 856
<< via3 >>
rect 6528 5982 6592 9406
rect 3138 5430 3279 5433
rect 3138 5368 3279 5430
rect 3138 5365 3279 5368
rect 651 4521 745 4658
rect 2483 4521 2577 4658
rect 1569 3474 1663 3611
rect -518 2018 -454 2218
rect 3714 2018 3778 2218
rect 1598 856 1662 1056
<< mimcap >>
rect 2880 9354 6280 9394
rect 2880 6034 2920 9354
rect 6240 6034 6280 9354
rect 2880 5994 6280 6034
<< mimcapcontact >>
rect 2920 6034 6240 9354
<< metal4 >>
rect 6512 9406 6608 9422
rect 2919 9354 6241 9355
rect 2919 6034 2920 9354
rect 6240 6034 6241 9354
rect 2919 6033 6241 6034
rect 3129 5434 3240 6033
rect 6512 5982 6528 9406
rect 6592 5982 6608 9406
rect 6512 5966 6608 5982
rect 3129 5433 3280 5434
rect 3129 5365 3138 5433
rect 3279 5430 3280 5433
rect 3279 5368 3348 5430
rect 3279 5365 3280 5368
rect 3129 5364 3280 5365
rect 374 4658 2578 4659
rect 374 4521 651 4658
rect 745 4521 2483 4658
rect 2577 4521 2578 4658
rect 374 4520 2578 4521
rect 374 3612 513 4520
rect 374 3611 1686 3612
rect 374 3474 1569 3611
rect 1663 3474 1686 3611
rect 374 3473 1686 3474
rect -519 2218 -453 2219
rect -519 2117 -518 2218
rect -971 2018 -518 2117
rect -454 2117 -453 2218
rect 374 2117 513 3473
rect 3713 2218 3779 2219
rect 3713 2117 3714 2218
rect -454 2018 3714 2117
rect 3778 2018 3779 2218
rect -971 2017 3779 2018
rect -971 955 -871 2017
rect 1597 1056 1663 1057
rect 1597 955 1598 1056
rect -971 856 1598 955
rect 1662 856 1663 1056
rect -971 855 1663 856
<< labels >>
rlabel metal2 4215 390 4215 390 3 vcc
port 1 e
rlabel metal2 463 6644 463 6644 7 vss
port 2 w
rlabel metal2 4778 4214 4778 4214 3 vo3
port 3 e
rlabel metal1 -66 4276 -66 4276 7 vd3
port 4 w
rlabel metal1 -66 4099 -66 4099 7 vd4
port 5 w
rlabel metal3 -66 4532 -66 4532 7 vb
port 6 w
rlabel metal3 2619 6975 2619 6975 7 vd1
port 7 w
<< end >>
