magic
tech sky130A
magscale 1 2
timestamp 1739144074
<< metal1 >>
rect 29697 5220 30542 5230
rect 29697 5130 30372 5220
rect 30362 4894 30372 5130
rect 30532 4894 30542 5220
<< via1 >>
rect 30372 4894 30532 5220
<< metal2 >>
rect 15595 9700 16395 9728
rect 10210 1481 10610 9697
rect 15595 9356 16020 9700
rect 16377 9356 16395 9700
rect 15595 9328 16395 9356
rect 29846 7166 30879 7176
rect 29846 6787 30097 7166
rect 29846 6777 30879 6787
rect 29846 6776 30246 6777
rect 30372 5220 30532 5230
rect 30372 4884 30532 4894
rect 14906 1993 15084 2336
rect 14906 1813 14944 1993
rect 15041 1813 15084 1993
rect 14906 1812 15084 1813
rect 14944 1803 15041 1812
rect 10210 1142 10251 1481
rect 10572 1142 10610 1481
rect 10210 1103 10610 1142
rect 13344 1493 21669 1503
rect 14082 1113 21669 1493
rect 13344 1104 21669 1113
rect 13344 1103 17814 1104
<< via2 >>
rect 16020 9356 16377 9700
rect 30097 6787 30879 7166
rect 30372 4894 30532 5220
rect 14944 1813 15041 1993
rect 10251 1142 10572 1481
rect 13344 1113 14082 1493
<< metal3 >>
rect 16010 9700 16387 9705
rect 16010 9356 16020 9700
rect 16377 9356 16387 9700
rect 16010 9351 16387 9356
rect 30087 6777 30097 7175
rect 30879 6777 30886 7175
rect 30362 5220 30542 5225
rect 30362 4894 30372 5220
rect 30532 4894 30542 5220
rect 30362 4889 30542 4894
rect 14934 1993 15051 1998
rect 14934 1813 14944 1993
rect 15041 1813 15051 1993
rect 14934 1808 15051 1813
rect 10241 1481 10582 1486
rect 10241 1142 10251 1481
rect 10572 1142 10582 1481
rect 10241 1137 10582 1142
rect 13334 1104 13344 1502
rect 14083 1104 14093 1502
rect 22607 1028 22787 1029
rect 18770 1027 22787 1028
rect 18770 849 18794 1027
rect 19276 849 22787 1027
rect 18770 848 22787 849
rect 23380 782 23560 1047
rect 23032 604 23042 782
rect 23524 604 23560 782
rect 23380 603 23560 604
rect 25838 782 26018 1032
rect 25838 604 25882 782
rect 26364 604 26374 782
rect 25838 603 26018 604
<< via3 >>
rect 16020 9356 16377 9700
rect 30097 7166 30879 7175
rect 30097 6787 30879 7166
rect 30097 6777 30879 6787
rect 30372 4894 30532 5220
rect 14944 1813 15041 1993
rect 10251 1142 10572 1481
rect 13344 1493 14083 1502
rect 13344 1113 14082 1493
rect 14082 1113 14083 1493
rect 13344 1104 14083 1113
rect 18794 849 19276 1027
rect 23042 604 23524 782
rect 25882 604 26364 782
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 14414 44152 14474 45152
rect 14966 44152 15026 45152
rect 15518 44152 15578 45152
rect 16070 44152 16130 45152
rect 16622 44152 16682 45152
rect 17174 44152 17234 45152
rect 17726 44152 17786 45152
rect 18278 44152 18338 45152
rect 18830 44152 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 400 43752 18890 44152
rect 400 1503 800 43752
rect 31400 9728 31800 44152
rect 15995 9700 31800 9728
rect 15995 9356 16020 9700
rect 16377 9356 31800 9700
rect 15995 9328 31800 9356
rect 31400 7176 31800 9328
rect 30005 7175 31800 7176
rect 30005 6777 30097 7175
rect 30879 6777 31800 7175
rect 30005 6776 31800 6777
rect 30362 5220 30542 5230
rect 30362 4894 30372 5220
rect 30532 4894 30542 5220
rect 14943 1993 15042 1994
rect 14943 1992 14944 1993
rect 14906 1813 14944 1992
rect 15041 1992 15042 1993
rect 15041 1813 15086 1992
rect 400 1502 14084 1503
rect 400 1481 13344 1502
rect 400 1142 10251 1481
rect 10572 1142 13344 1481
rect 400 1104 13344 1142
rect 14083 1104 14084 1502
rect 400 1103 14084 1104
rect 400 1000 800 1103
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 1813
rect 18770 1027 19277 1028
rect 18770 849 18794 1027
rect 19276 849 19277 1027
rect 18770 848 19277 849
rect 18770 0 18950 848
rect 22634 782 23560 783
rect 22634 604 23042 782
rect 23524 604 23560 782
rect 22634 603 23560 604
rect 25838 782 26678 783
rect 25838 604 25882 782
rect 26364 604 26678 782
rect 25838 603 26678 604
rect 22634 0 22814 603
rect 26498 0 26678 603
rect 30362 0 30542 4894
rect 31400 1000 31800 6776
use BGR_BJT_final  BGR_BJT_final_0 ~/Dalin/gds_files/tinytape_diff_BGR/tt_um_DalinEM_diff_amp/mag/BGR_BJT_final
timestamp 1739140642
transform 0 -1 16030 -1 0 9692
box -168 -2 7713 5682
use diff_final_v0  diff_final_v0_0 ~/Dalin/Projects/tinytape/diff_files
timestamp 1738105933
transform 1 0 10675 0 1 3795
box 10993 -2832 19171 3381
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 31400 1000 31800 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 1000 800 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
