** sch_path: /home/zerotoasic/Dalin/Projects/tinytape/voltage_ref_BJT/BGR_BJT_stage2.sch
.subckt BGR_BJT_stage2 vcc vr vref vref0 vss
*.PININFO vref:O vcc:I vss:I vref0:I vr:I
XM4 net2 net3 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM5 net3 net3 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM6 net1 net4 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM7 net4 net4 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM10 net3 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM11 net4 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM12 vref vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM16 net5 net6 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM15 net6 net6 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM14 net6 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM19 vref net7 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM18 net7 net7 vref vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM17 net7 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM1 net3 net3 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM2 net3 net3 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM3 net3 net3 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM8 net4 net4 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM9 net4 net4 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM13 net4 net4 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM20 net6 net6 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM21 net6 net6 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM22 net6 net6 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM23 net7 net7 vref vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM24 net7 net7 vref vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM25 net7 net7 vref vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
.ends
.end
