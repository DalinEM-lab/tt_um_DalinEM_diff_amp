* NGSPICE file created from tt_um_DalinEM_diff_amp.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_58FN7G a_n1800_n277# a_1800_n180# a_n1858_n180#
+ w_n1894_n280#
X0 a_1800_n180# a_n1800_n277# a_n1858_n180# w_n1894_n280# sky130_fd_pr__pfet_01v8_lvt ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=18
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_59CFV9 a_1200_n600# a_n1258_n600# a_n1200_n688#
+ VSUBS
X0 a_1200_n600# a_n1200_n688# a_n1258_n600# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=12
.ends

.subckt sky130_fd_pr__nfet_01v8_Q93DRV a_n558_n300# a_n500_n388# a_n660_n474# a_500_n300#
X0 a_500_n300# a_n500_n388# a_n558_n300# a_n660_n474# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=5
.ends

.subckt diff_final_v0 vout vin_p vin_n vb vcc vss
Xsky130_fd_pr__pfet_01v8_lvt_58FN7G_0 m1_15336_1751# vout vcc vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM1 m1_11317_n793# m1_15336_1751# vin_p vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM2 m1_11317_n793# vout vin_n vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM3 vss vb vss m1_11317_n793# sky130_fd_pr__nfet_01v8_Q93DRV
XXM4 m1_15336_1751# vcc vout vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM5 m1_15336_1751# vcc m1_15336_1751# vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM6 m1_15336_1751# m1_15336_1751# vcc vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
Xsky130_fd_pr__nfet_01v8_lvt_59CFV9_0 vout m1_11317_n793# vin_n vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM8 m1_15336_1751# m1_11317_n793# vin_p vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
.ends

.subckt tt_um_DalinEM_diff_amp clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] VDPWR VGND
Xdiff_final_v0_0 ua[0] ua[1] ua[2] ua[3] VDPWR VGND diff_final_v0
.ends

