magic
tech sky130A
magscale 1 2
timestamp 1740710330
<< locali >>
rect 2075 2434 6860 2445
rect 2049 1894 6860 2434
rect 2075 1889 6860 1894
<< metal1 >>
rect 2168 779 2431 825
<< metal2 >>
rect 102 5372 161 5566
rect 1842 2246 1922 2256
rect 1842 1523 1922 2162
rect 1842 1443 2041 1523
rect 7692 965 7710 1014
rect 83 22 139 186
rect 2134 130 2478 290
<< via2 >>
rect 1842 2162 1922 2246
<< metal3 >>
rect 1832 2246 1932 2251
rect 1546 2162 1842 2246
rect 1922 2162 1932 2246
rect 1832 2157 1932 2162
use BGR_BJT_stage1  BGR_BJT_stage1_0 ~/Project_tinytape/magic/mag/BGR_BJT_final/layout_BGR_BJT_stage1
timestamp 1739137757
transform 1 0 -5377 0 1 3366
box 5349 -3380 12358 2268
use BGR_BJT_stage2  BGR_BJT_stage2_0 ~/Project_tinytape/magic/mag/BGR_BJT_final/layout_BGR_BJT_stage-2
timestamp 1739131682
transform 1 0 2947 0 -1 2436
box -928 535 4746 2353
<< labels >>
rlabel metal2 85 102 85 102 7 vcc
port 1 w
rlabel metal2 103 5468 103 5468 7 vss
port 2 w
rlabel metal2 7709 990 7709 990 7 vref
port 3 w
<< end >>
