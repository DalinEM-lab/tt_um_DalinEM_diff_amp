magic
tech sky130A
magscale 1 2
timestamp 1741224555
<< nwell >>
rect 6472 -3262 9085 4497
<< psubdiff >>
rect 6617 -3656 6677 -3622
rect 14846 -3656 14906 -3622
rect 6617 -3682 6651 -3656
rect 6617 -4931 6651 -4905
rect 14872 -3682 14906 -3656
rect 14872 -4931 14906 -4905
rect 6617 -4965 6677 -4931
rect 14846 -4965 14906 -4931
<< nsubdiff >>
rect 6565 4397 6625 4431
rect 8905 4397 8965 4431
rect 6565 4371 6599 4397
rect 6565 -3190 6599 -3164
rect 8931 4371 8965 4397
rect 8931 -3190 8965 -3164
rect 6565 -3224 6625 -3190
rect 8905 -3224 8965 -3190
<< psubdiffcont >>
rect 6677 -3656 14846 -3622
rect 6617 -4905 6651 -3682
rect 14872 -4905 14906 -3682
rect 6677 -4965 14846 -4931
<< nsubdiffcont >>
rect 6625 4397 8905 4431
rect 6565 -3164 6599 4371
rect 8931 -3164 8965 4371
rect 6625 -3224 8905 -3190
<< locali >>
rect 6457 4501 9122 4514
rect 6457 890 6491 4501
rect 9083 4298 9122 4501
rect 6656 4280 8931 4298
rect 6656 890 6691 4280
rect 6457 72 6565 890
rect 6599 72 6691 890
rect 6457 -3104 6508 72
rect 6457 -3280 6507 -3104
rect 6656 -3123 6691 72
rect 8806 3719 8931 4280
rect 8965 3719 9122 4298
rect 8806 1239 8871 3719
rect 9013 1239 9122 3719
rect 8806 -514 8931 1239
rect 8965 -514 9122 1239
rect 8806 -2994 8887 -514
rect 9029 -925 9122 -514
rect 9029 -1012 13862 -925
rect 13819 -1013 13862 -1012
rect 9029 -1391 11291 -1304
rect 9029 -2994 9122 -1391
rect 8806 -3123 8931 -2994
rect 6656 -3137 8931 -3123
rect 8965 -3137 9122 -2994
rect 9072 -3261 9122 -3137
rect 6457 -3281 6620 -3280
rect 9072 -3281 9108 -3261
rect 6457 -3288 9108 -3281
rect 11246 -3294 11291 -1391
rect 11524 -1391 13542 -1304
rect 11524 -3034 11588 -1391
rect 13428 -2820 13542 -1391
rect 13829 -2820 13862 -1013
rect 13428 -3034 13862 -2820
rect 11524 -3054 13862 -3034
rect 11524 -3060 13866 -3054
rect 11246 -3296 11376 -3294
rect 13439 -3296 13866 -3060
rect 11246 -3310 13866 -3296
rect 6553 -3619 14389 -3582
rect 6553 -5119 6563 -3619
rect 6710 -3622 14389 -3619
rect 14505 -3622 14960 -3582
rect 14846 -3656 14960 -3622
rect 14505 -3682 14960 -3656
rect 6710 -3743 14389 -3731
rect 14505 -3743 14872 -3682
rect 6710 -3769 14872 -3743
rect 6710 -4847 6731 -3769
rect 14791 -4847 14872 -3769
rect 6710 -4905 14872 -4847
rect 14906 -4905 14960 -3682
rect 6710 -4921 14960 -4905
rect 6804 -4922 14960 -4921
rect 14482 -4931 14960 -4922
rect 14846 -4965 14960 -4931
rect 14482 -5119 14960 -4965
rect 6553 -5136 14960 -5119
rect 6562 -5137 14960 -5136
<< viali >>
rect 6491 4431 9083 4501
rect 6491 4397 6625 4431
rect 6625 4397 8905 4431
rect 8905 4397 9083 4431
rect 6491 4371 9083 4397
rect 6491 890 6565 4371
rect 6565 890 6599 4371
rect 6599 4298 8931 4371
rect 8931 4298 8965 4371
rect 8965 4298 9083 4371
rect 6599 890 6656 4298
rect 6508 -3104 6565 72
rect 6507 -3164 6565 -3104
rect 6565 -3164 6599 72
rect 6599 -3137 6656 72
rect 8871 1239 8931 3719
rect 8931 1239 8965 3719
rect 8965 1239 9013 3719
rect 8887 -2994 8931 -514
rect 8931 -2994 8965 -514
rect 8965 -1012 9029 -514
rect 8965 -1013 13819 -1012
rect 8965 -1304 13829 -1013
rect 8965 -2994 9029 -1304
rect 6599 -3164 8931 -3137
rect 8931 -3164 8965 -3137
rect 8965 -3164 9072 -3137
rect 6507 -3190 9072 -3164
rect 6507 -3224 6625 -3190
rect 6625 -3224 8905 -3190
rect 8905 -3224 9072 -3190
rect 6507 -3280 9072 -3224
rect 6620 -3281 9072 -3280
rect 11291 -3060 11524 -1304
rect 13542 -2820 13829 -1304
rect 11291 -3294 13439 -3060
rect 11376 -3296 13439 -3294
rect 6563 -3622 6710 -3619
rect 14389 -3622 14505 -3582
rect 6563 -3656 6677 -3622
rect 6677 -3627 6710 -3622
rect 6677 -3628 6839 -3627
rect 14389 -3628 14505 -3622
rect 6677 -3656 14505 -3628
rect 6563 -3682 14505 -3656
rect 6563 -4905 6617 -3682
rect 6617 -4905 6651 -3682
rect 6651 -3731 14505 -3682
rect 6651 -4905 6710 -3731
rect 14389 -3743 14505 -3731
rect 6563 -4921 6710 -4905
rect 6563 -4922 6804 -4921
rect 6563 -4931 14482 -4922
rect 6563 -4965 6677 -4931
rect 6677 -4965 14482 -4931
rect 6563 -5119 14482 -4965
<< metal1 >>
rect 6479 4501 9095 4507
rect 6479 4292 6491 4501
rect 9083 4298 9095 4501
rect 6481 890 6491 4292
rect 6656 4292 9095 4298
rect 6656 890 6666 4292
rect 6803 1029 6813 2029
rect 6877 1029 6887 2029
rect 6951 979 7156 4069
rect 7238 3405 7248 4005
rect 7320 3405 7330 4005
rect 7404 979 7609 4069
rect 7680 2266 7690 3266
rect 7754 2266 7764 3266
rect 7840 979 8045 4069
rect 8114 3405 8124 4005
rect 8196 3405 8206 4005
rect 8280 979 8485 4064
rect 8865 3719 9019 3731
rect 8556 1029 8566 2029
rect 8630 1029 8640 2029
rect 8865 1239 8871 3719
rect 9013 1239 9019 3719
rect 8865 1227 9019 1239
rect 6881 927 6891 979
rect 7171 927 7181 979
rect 7319 927 7329 979
rect 7609 927 7619 979
rect 7757 927 7767 979
rect 8047 927 8057 979
rect 8195 927 8205 979
rect 8485 927 8495 979
rect 6485 878 6662 890
rect 6296 634 6891 734
rect 6991 634 7577 734
rect 7677 634 8015 734
rect 8115 634 8205 734
rect 8305 634 10030 734
rect 10312 634 10322 734
rect 6296 325 7139 425
rect 7239 325 7329 425
rect 7429 325 7767 425
rect 7867 325 8453 425
rect 8553 325 8710 425
rect 6502 72 6662 84
rect 6949 78 6959 130
rect 7239 78 7249 130
rect 7387 78 7397 130
rect 7677 78 7687 130
rect 7825 78 7835 130
rect 8115 78 8125 130
rect 8263 78 8273 130
rect 8553 78 8563 130
rect 6498 -3104 6508 72
rect 6497 -3280 6507 -3104
rect 6656 -3131 6666 72
rect 6804 -972 6814 28
rect 6878 -972 6888 28
rect 6955 -3004 7160 78
rect 7238 -2948 7248 -2348
rect 7320 -2948 7330 -2348
rect 7408 -3004 7613 78
rect 7680 -2132 7690 -1132
rect 7754 -2132 7764 -1132
rect 7844 -3008 8049 78
rect 8113 -2948 8123 -2348
rect 8195 -2948 8205 -2348
rect 8276 -3004 8481 78
rect 8556 -972 8566 28
rect 8630 -972 8640 28
rect 8881 -514 9035 -502
rect 8881 -2994 8887 -514
rect 9029 -1006 9035 -514
rect 13536 -1006 13835 -1001
rect 9029 -1012 13835 -1006
rect 13819 -1013 13835 -1012
rect 9029 -1310 11291 -1304
rect 9029 -2994 9035 -1310
rect 8881 -3006 9035 -2994
rect 6656 -3137 9084 -3131
rect 6501 -3281 6620 -3280
rect 9072 -3281 9084 -3137
rect 6501 -3287 9084 -3281
rect 6501 -3292 6662 -3287
rect 11285 -3294 11291 -1310
rect 11524 -1310 13542 -1304
rect 11524 -3054 11530 -1310
rect 11639 -2526 11649 -1526
rect 11701 -2526 11711 -1526
rect 11776 -2961 11977 -1461
rect 12057 -2902 12067 -1902
rect 12119 -2902 12129 -1902
rect 12053 -3001 12134 -2955
rect 12195 -2970 12396 -1470
rect 12475 -2526 12485 -1526
rect 12537 -2526 12547 -1526
rect 12475 -3001 12556 -2955
rect 12618 -2966 12819 -1466
rect 12893 -2902 12903 -1902
rect 12955 -2902 12965 -1902
rect 12888 -3001 12969 -2955
rect 13024 -2966 13225 -1466
rect 13311 -2526 13321 -1526
rect 13373 -2526 13383 -1526
rect 13532 -2820 13542 -1310
rect 13829 -2820 13839 -1013
rect 13536 -2832 13835 -2820
rect 13519 -2955 13529 -2946
rect 13266 -3001 13529 -2955
rect 13519 -3005 13529 -3001
rect 13653 -3005 13663 -2946
rect 11524 -3060 13451 -3054
rect 11285 -3296 11376 -3294
rect 13439 -3296 13451 -3060
rect 11285 -3302 13451 -3296
rect 11285 -3306 11530 -3302
rect 14383 -3582 14511 -3563
rect 6557 -3619 6716 -3607
rect 6553 -4915 6563 -3619
rect 6710 -3621 6720 -3619
rect 6710 -3622 6851 -3621
rect 14373 -3622 14383 -3582
rect 6710 -3627 14383 -3622
rect 6839 -3628 14383 -3627
rect 6551 -5119 6563 -4915
rect 6710 -3737 14383 -3731
rect 6710 -4915 6720 -3737
rect 14373 -3765 14383 -3737
rect 14530 -3765 14540 -3582
rect 6814 -4098 6824 -3998
rect 6888 -4098 6898 -3998
rect 7109 -4325 8528 -3944
rect 8758 -4098 8768 -3998
rect 8820 -4098 8830 -3998
rect 6814 -4684 6824 -4584
rect 6888 -4684 6898 -4584
rect 6833 -4728 6879 -4694
rect 6833 -4774 6911 -4728
rect 7113 -4739 8532 -4358
rect 8759 -4364 8838 -4318
rect 9143 -4325 10562 -3944
rect 10688 -3954 10781 -3908
rect 10709 -3994 10755 -3954
rect 10690 -4274 10700 -4174
rect 10764 -4274 10774 -4174
rect 8758 -4684 8768 -4584
rect 8820 -4684 8830 -4584
rect 9139 -4735 10558 -4354
rect 10697 -4364 10776 -4318
rect 10972 -4320 12391 -3939
rect 12634 -4098 12644 -3998
rect 12696 -4098 12706 -3998
rect 10690 -4508 10700 -4408
rect 10764 -4508 10774 -4408
rect 10972 -4735 12391 -4354
rect 12636 -4364 12715 -4318
rect 12942 -4325 14361 -3944
rect 14566 -4098 14576 -3998
rect 14640 -4098 14650 -3998
rect 12634 -4684 12644 -4584
rect 12696 -4684 12706 -4584
rect 12942 -4731 14361 -4350
rect 14566 -4684 14576 -4584
rect 14640 -4684 14650 -4584
rect 14585 -4728 14631 -4691
rect 14552 -4774 14631 -4728
rect 6710 -4916 6816 -4915
rect 6710 -4921 14494 -4916
rect 6804 -4922 14494 -4921
rect 14482 -5119 14494 -4922
rect 6551 -5125 14494 -5119
<< via1 >>
rect 6491 4298 9083 4501
rect 6491 890 6656 4298
rect 6813 1029 6877 2029
rect 7248 3405 7320 4005
rect 7690 2266 7754 3266
rect 8124 3405 8196 4005
rect 8566 1029 8630 2029
rect 6891 927 7171 979
rect 7329 927 7609 979
rect 7767 927 8047 979
rect 8205 927 8485 979
rect 6891 634 6991 734
rect 7577 634 7677 734
rect 8015 634 8115 734
rect 8205 634 8305 734
rect 10030 634 10312 734
rect 7139 325 7239 425
rect 7329 325 7429 425
rect 7767 325 7867 425
rect 8453 325 8553 425
rect 6959 78 7239 130
rect 7397 78 7677 130
rect 7835 78 8115 130
rect 8273 78 8553 130
rect 6508 -3104 6656 72
rect 6507 -3137 6656 -3104
rect 6814 -972 6878 28
rect 7248 -2948 7320 -2348
rect 7690 -2132 7754 -1132
rect 8123 -2948 8195 -2348
rect 8566 -972 8630 28
rect 10166 -1304 13829 -1013
rect 6507 -3280 9072 -3137
rect 6620 -3281 9072 -3280
rect 11649 -2526 11701 -1526
rect 12067 -2902 12119 -1902
rect 12485 -2526 12537 -1526
rect 12903 -2902 12955 -1902
rect 13321 -2526 13373 -1526
rect 13542 -2820 13829 -1304
rect 13529 -3005 13653 -2946
rect 11376 -3296 13439 -3060
rect 6563 -3627 6710 -3619
rect 6563 -3628 6839 -3627
rect 14383 -3628 14389 -3582
rect 14389 -3628 14505 -3582
rect 6563 -3731 14505 -3628
rect 6563 -4921 6710 -3731
rect 14383 -3743 14389 -3731
rect 14389 -3743 14505 -3731
rect 14505 -3743 14530 -3582
rect 14383 -3765 14530 -3743
rect 6824 -4098 6888 -3998
rect 8768 -4098 8820 -3998
rect 6824 -4684 6888 -4584
rect 10700 -4274 10764 -4174
rect 8768 -4684 8820 -4584
rect 12644 -4098 12696 -3998
rect 10700 -4508 10764 -4408
rect 14576 -4098 14640 -3998
rect 12644 -4684 12696 -4584
rect 14576 -4684 14640 -4584
rect 6563 -4922 6804 -4921
rect 6563 -5119 14482 -4922
<< metal2 >>
rect 6402 4501 9083 4511
rect 6402 4287 6491 4501
rect 6656 4288 9083 4298
rect 7248 4005 9929 4015
rect 7320 3915 8124 4005
rect 7248 3395 7320 3405
rect 8196 3915 9929 4005
rect 8124 3395 8196 3405
rect 7690 3266 7754 3276
rect 7690 2256 7754 2266
rect 6813 2029 6877 2039
rect 6813 1019 6877 1029
rect 8566 2029 8630 2039
rect 8566 1019 8630 1029
rect 6491 880 6656 890
rect 6891 979 7171 989
rect 6891 917 7171 927
rect 7329 979 7609 989
rect 7329 917 7609 927
rect 7767 979 8047 989
rect 7767 917 8047 927
rect 8205 979 8485 989
rect 8205 917 8485 927
rect 6891 734 6991 917
rect 6891 624 6991 634
rect 7139 425 7239 435
rect 7139 140 7239 325
rect 7329 425 7429 917
rect 7329 315 7429 325
rect 7577 734 7677 744
rect 7577 140 7677 634
rect 7767 425 7867 917
rect 7767 315 7867 325
rect 8015 734 8115 744
rect 8015 140 8115 634
rect 8205 734 8305 917
rect 8205 624 8305 634
rect 8453 425 8553 435
rect 8453 140 8553 325
rect 6959 130 7239 140
rect 6508 72 6656 82
rect 6507 -3104 6508 -3094
rect 6959 68 7239 78
rect 7397 130 7677 140
rect 7397 68 7677 78
rect 7835 130 8115 140
rect 7835 68 8115 78
rect 8273 130 8553 140
rect 8273 68 8553 78
rect 6814 28 6878 38
rect 6814 -982 6878 -972
rect 8566 28 8630 38
rect 8566 -982 8630 -972
rect 7690 -1132 7754 -1122
rect 7690 -2142 7754 -2132
rect 9829 -1516 9929 3915
rect 10020 734 10312 744
rect 10020 624 10312 634
rect 10166 -1013 13829 -1003
rect 10166 -1314 13542 -1304
rect 9829 -1526 13373 -1516
rect 9829 -1616 11649 -1526
rect 7248 -2338 8648 -2337
rect 9829 -2338 9929 -1616
rect 7248 -2348 9929 -2338
rect 7320 -2437 8123 -2348
rect 7248 -2958 7320 -2948
rect 8195 -2437 9929 -2348
rect 8520 -2438 9929 -2437
rect 11701 -1616 12485 -1526
rect 11649 -2536 11701 -2526
rect 12067 -1902 12119 -1892
rect 8123 -2958 8195 -2948
rect 12537 -1616 13321 -1526
rect 12485 -2536 12537 -2526
rect 12903 -1902 12955 -1892
rect 12067 -3050 12119 -2902
rect 13321 -2536 13373 -2526
rect 13542 -2830 13829 -2820
rect 12903 -3050 12955 -2902
rect 13529 -2946 15141 -2936
rect 13653 -3005 15141 -2946
rect 13529 -3015 15141 -3005
rect 11376 -3060 13439 -3050
rect 6656 -3137 9072 -3127
rect 6507 -3281 6620 -3280
rect 6507 -3290 9072 -3281
rect 6620 -3291 9072 -3290
rect 11376 -3306 13439 -3296
rect 14383 -3582 14530 -3572
rect 6563 -3617 6710 -3609
rect 6563 -3618 6839 -3617
rect 6563 -3619 14383 -3618
rect 6710 -3627 14383 -3619
rect 6839 -3628 14383 -3627
rect 6497 -5119 6563 -4911
rect 6710 -3741 14383 -3731
rect 6824 -3998 6888 -3988
rect 6824 -4108 6888 -4098
rect 8768 -3998 8820 -3741
rect 8768 -4108 8820 -4098
rect 12644 -3998 12696 -3741
rect 14383 -3775 14530 -3765
rect 12644 -4108 12696 -4098
rect 14576 -3998 14640 -3988
rect 14576 -4108 14640 -4098
rect 10700 -4174 10764 -4164
rect 10700 -4284 10764 -4274
rect 10700 -4408 10764 -4398
rect 10700 -4518 10764 -4508
rect 6824 -4584 6888 -4574
rect 6824 -4694 6888 -4684
rect 8768 -4584 8820 -4574
rect 6710 -4912 6804 -4911
rect 8768 -4912 8820 -4684
rect 12644 -4584 12696 -4574
rect 12644 -4912 12696 -4684
rect 14576 -4584 14640 -4574
rect 14576 -4694 14640 -4684
rect 6710 -4921 14482 -4912
rect 6804 -4922 14482 -4921
rect 15062 -5083 15141 -3015
rect 6497 -5129 14482 -5119
<< via2 >>
rect 7690 2266 7754 3266
rect 6813 1029 6877 2029
rect 8566 1029 8630 2029
rect 6814 -972 6878 28
rect 8566 -972 8630 28
rect 7690 -2132 7754 -1132
rect 10020 634 10030 734
rect 10030 634 10312 734
rect 6824 -4098 6888 -3998
rect 14576 -4098 14640 -3998
rect 10700 -4274 10764 -4174
rect 10700 -4508 10764 -4408
rect 6824 -4684 6888 -4584
rect 14576 -4684 14640 -4584
<< metal3 >>
rect 7680 3266 7764 3271
rect 7680 2266 7690 3266
rect 7754 2352 7764 3266
rect 7754 2266 8872 2352
rect 7680 2261 8872 2266
rect 7694 2252 8872 2261
rect 6803 2029 6887 2034
rect 6803 1029 6813 2029
rect 6877 1029 6887 2029
rect 6803 1024 6887 1029
rect 8556 2029 8640 2034
rect 8556 1029 8566 2029
rect 8630 1029 8640 2029
rect 8556 1024 8640 1029
rect 8772 36 8872 2252
rect 10010 734 11270 739
rect 10010 634 10020 734
rect 10312 634 11270 734
rect 10010 629 11270 634
rect 8772 33 8963 36
rect 6804 28 8963 33
rect 6804 -972 6814 28
rect 6878 -67 8566 28
rect 6878 -972 6888 -67
rect 6804 -977 6888 -972
rect 8556 -972 8566 -67
rect 8630 -67 8963 28
rect 8630 -972 8640 -67
rect 8556 -977 8640 -972
rect 7680 -1132 7764 -1127
rect 7680 -2132 7690 -1132
rect 7754 -2132 7764 -1132
rect 7680 -2137 7764 -2132
rect 6807 -3998 6905 -3993
rect 6807 -4098 6824 -3998
rect 6888 -4098 6905 -3998
rect 6807 -4103 6905 -4098
rect 8853 -4169 8963 -67
rect 14538 -3998 14666 -3993
rect 14538 -4098 14576 -3998
rect 14640 -4098 14666 -3998
rect 14538 -4103 14666 -4098
rect 8853 -4174 15036 -4169
rect 8853 -4274 10700 -4174
rect 10764 -4274 15036 -4174
rect 8853 -4279 15036 -4274
rect 14926 -4355 15036 -4279
rect 10674 -4408 10789 -4403
rect 10674 -4508 10700 -4408
rect 10764 -4508 10789 -4408
rect 10674 -4513 10789 -4508
rect 14926 -4455 15454 -4355
rect 14926 -4579 15036 -4455
rect 6814 -4584 15036 -4579
rect 6814 -4684 6824 -4584
rect 6888 -4684 14576 -4584
rect 14640 -4684 15036 -4584
rect 6814 -4689 15036 -4684
<< via3 >>
rect 6813 1029 6877 2029
rect 8566 1029 8630 2029
rect 7690 -2132 7754 -1132
rect 6824 -4098 6888 -3998
rect 14576 -4098 14640 -3998
rect 10700 -4508 10764 -4408
<< metal4 >>
rect 6812 2029 6878 2030
rect 6812 1029 6813 2029
rect 6877 1128 6878 2029
rect 8565 2029 8631 2030
rect 8565 1128 8566 2029
rect 6877 1029 8566 1128
rect 8630 1128 8631 2029
rect 8630 1029 9266 1128
rect 6812 1028 9266 1029
rect 7689 -1132 7755 -1131
rect 7689 -2132 7690 -1132
rect 7754 -1166 7755 -1132
rect 9166 -1166 9266 1028
rect 13250 533 14658 599
rect 7754 -1266 9266 -1166
rect 14592 -1180 14658 533
rect 7754 -2132 7755 -1266
rect 7689 -2133 7755 -2132
rect 9166 -3997 9266 -1266
rect 14591 -1258 14658 -1180
rect 14591 -3997 14657 -1258
rect 6823 -3998 15304 -3997
rect 6823 -4098 6824 -3998
rect 6888 -4098 14576 -3998
rect 14640 -4098 15304 -3998
rect 6823 -4099 15304 -4098
rect 15202 -4169 15304 -4099
rect 15202 -4269 15454 -4169
rect 15202 -4407 15304 -4269
rect 10699 -4408 15304 -4407
rect 10699 -4508 10700 -4408
rect 10764 -4508 15304 -4408
rect 10699 -4509 15304 -4508
use sky130_fd_pr__nfet_01v8_lvt_AR4WA2  sky130_fd_pr__nfet_01v8_lvt_AR4WA2_0
timestamp 1740448279
transform 1 0 13639 0 1 -4136
box -998 -238 998 238
use sky130_fd_pr__pfet_01v8_lvt_NH7ZMU  sky130_fd_pr__pfet_01v8_lvt_NH7ZMU_0
timestamp 1740449209
transform 1 0 7941 0 1 -1460
box -284 -1600 284 1600
use sky130_fd_pr__pfet_01v8_lvt_NH7ZMU  sky130_fd_pr__pfet_01v8_lvt_NH7ZMU_1
timestamp 1740449209
transform 1 0 8379 0 1 2517
box -284 -1600 284 1600
use sky130_fd_pr__cap_mim_m3_1_FGZHLY  XC1
timestamp 1741206728
transform 0 -1 12295 1 0 1601
box -1186 -1040 1186 1040
use sky130_fd_pr__pfet_01v8_6JHA76  XM3
timestamp 1740447052
transform 1 0 12511 0 1 -2214
box -1003 -919 1003 919
use sky130_fd_pr__pfet_01v8_lvt_NH7ZMU  XM4
timestamp 1740449209
transform 1 0 7503 0 1 2517
box -284 -1600 284 1600
use sky130_fd_pr__pfet_01v8_lvt_NH7ZMU  XM5
timestamp 1740449209
transform 1 0 7941 0 1 2517
box -284 -1600 284 1600
use sky130_fd_pr__pfet_01v8_lvt_NH7ZMU  XM7
timestamp 1740449209
transform 1 0 7065 0 1 -1460
box -284 -1600 284 1600
use sky130_fd_pr__pfet_01v8_lvt_NH7ZMU  XM8
timestamp 1740449209
transform 1 0 7065 0 1 2517
box -284 -1600 284 1600
use sky130_fd_pr__nfet_01v8_lvt_AR4WA2  XM9
timestamp 1740448279
transform 1 0 7825 0 1 -4546
box -998 -238 998 238
use sky130_fd_pr__nfet_01v8_lvt_AR4WA2  XM10
timestamp 1740448279
transform 1 0 9763 0 1 -4546
box -998 -238 998 238
use sky130_fd_pr__pfet_01v8_lvt_NH7ZMU  XM11
timestamp 1740449209
transform 1 0 8379 0 1 -1460
box -284 -1600 284 1600
use sky130_fd_pr__pfet_01v8_lvt_NH7ZMU  XM12
timestamp 1740449209
transform 1 0 7503 0 1 -1460
box -284 -1600 284 1600
use sky130_fd_pr__nfet_01v8_lvt_AR4WA2  XM15
timestamp 1740448279
transform 1 0 13639 0 1 -4546
box -998 -238 998 238
use sky130_fd_pr__nfet_01v8_lvt_AR4WA2  XM16
timestamp 1740448279
transform 1 0 9763 0 1 -4136
box -998 -238 998 238
use sky130_fd_pr__nfet_01v8_lvt_AR4WA2  XM17
timestamp 1740448279
transform 1 0 11701 0 1 -4136
box -998 -238 998 238
use sky130_fd_pr__nfet_01v8_lvt_AR4WA2  XM18
timestamp 1740448279
transform 1 0 11701 0 1 -4546
box -998 -238 998 238
use sky130_fd_pr__nfet_01v8_lvt_AR4WA2  XM19
timestamp 1740448279
transform 1 0 7825 0 1 -4136
box -998 -238 998 238
<< labels >>
rlabel metal2 6403 4400 6403 4400 7 vcc
port 1 w
rlabel metal2 6499 -5026 6499 -5026 7 vss
port 2 w
rlabel metal1 6298 686 6298 686 7 vd1
port 3 w
rlabel metal1 6297 371 6297 371 7 vd2
port 4 w
rlabel metal4 15453 -4218 15453 -4218 7 vd4
port 5 w
rlabel metal3 15452 -4406 15452 -4406 7 vd3
port 6 w
rlabel metal2 15098 -5081 15098 -5081 5 vb1
port 7 s
<< end >>
