* NGSPICE file created from tt_um_DalinEM_test_flat.ext - technology: sky130A

.subckt tt_um_DalinEM_test_flat ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] VDPWR VGND
X0 3_OTA_0.3rd_3_OTA_0.vd3.t9 3_OTA_0.3rd_3_OTA_0.vd3.t8 VGND.t80 VGND.t73 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X1 a_18163_10306.t4 ua[2].t0 a_18046_7223# VGND.t13 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X2 VGND.t86 a_12378_15906.t38 a_12378_15906.t39 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t32 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t5 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X4 3_OTA_0.OTA_vref_0.vb 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t20 VDPWR.t63 VDPWR.t51 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X5 a_24889_22946.t1 3_OTA_0.OTA_stage1_0.vd1 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X6 a_12378_15906.t43 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t16 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X7 a_3013_4521.t44 a_3013_4521.t43 VGND.t53 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X8 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t29 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 a_3013_4521.t10 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X9 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t31 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t18 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X10 a_3013_4521.t42 a_3013_4521.t41 VGND.t44 VGND.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X11 a_12564_25551.t11 3_OTA_0.OTA_vref_0.vb1.t6 VDPWR.t45 VDPWR.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=81200,2916
X12 a_12564_25551.t5 3_OTA_0.OTA_stage1_0.vd1.t0 3_OTA_0.3rd_3_OTA_0.vd4.t3 VDPWR.t37 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X13 a_12378_15906.t47 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t15 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X14 a_6719_5623# a_6631_5681# a_6631_5681# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X15 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t28 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 a_3013_4521.t12 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X16 a_15996_17227# 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t21 VDPWR.t62 VDPWR.t61 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X17 VGND.t36 a_3013_4521.t39 a_3013_4521.t40 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X18 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t0 a_6631_6971# a_6719_6913# VGND.t26 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=11600,516
X19 3_OTA_0.OTA_stage1_0.vd1 3_OTA_0.OTA_stage1_0.vd2.t0 VDPWR.t24 VDPWR.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X20 ua[1].t1 a_18163_10306.t0 VDPWR.t36 VDPWR.t34 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X21 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t27 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 a_3013_4521.t11 VGND.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X22 a_15996_21097# a_15996_21097# 3_OTA_0.OTA_vref_0.vb VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=5800,258 d=5800,258
X23 a_16084_17427# a_15996_17227# a_15996_17227# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X24 a_12378_15906.t37 a_12378_15906.t36 VGND.t46 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X25 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t12 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t15 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X26 a_24889_22946.t0 ua[0].t1 VGND.t40 sky130_fd_pr__res_xhigh_po_0p35 l=1.2
X27 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t6 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t30 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X28 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t26 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 a_3013_4521.t6 VGND.t19 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X29 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t25 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 a_3013_4521.t7 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X30 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t29 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t16 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X31 ua[1].t3 ua[3].t0 a_18046_7223# VGND.t48 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X32 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t14 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t28 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X33 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t22 VDPWR.t60 VDPWR.t59 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=11600,516
X34 VGND.t79 3_OTA_0.3rd_3_OTA_0.vd3.t12 3_OTA_0.3rd_3_OTA_0.vd4.t7 VGND.t71 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X35 VDPWR.t9 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t20 a_6631_6971# VDPWR.t8 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X36 3_OTA_0.3rd_3_OTA_0.vd3.t0 3_OTA_0.OTA_stage1_0.vd2.t4 a_12564_25551.t0 VDPWR.t38 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X37 VDPWR.t1 a_21048_25880.t10 a_21048_25880.t11 VDPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X38 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t14 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 a_12378_15906.t0 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X39 a_6719_4333# a_6631_4391# a_6631_4391# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X40 a_18163_10306.t1 a_18163_10306.t0 VDPWR.t35 VDPWR.t34 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X41 3_OTA_0.OTA_stage1_0.vd2.t3 3_OTA_0.OTA_stage1_0.vd2.t0 VDPWR.t23 VDPWR.t22 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X42 a_12378_15906.t35 a_12378_15906.t34 VGND.t4 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X43 VDPWR.t7 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t21 a_6631_4391# VDPWR.t6 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X44 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t5 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t14 VGND.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X45 a_6631_5681# a_6631_5681# a_6719_5623# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X46 a_3013_4521.t5 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t24 VGND.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X47 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t10 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t13 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X48 VGND.t60 3_OTA_0.OTA_vref_0.vb a_22654_21988# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=1.048143 ps=7.775429 w=5.5 l=1.5
**devattr s=63800,2316 d=31900,1158
X49 3_OTA_0.OTA_stage1_0.vd1 ua[3].t1 a_3537_27009# VGND.t30 sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.58 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X50 a_22654_21988# 3_OTA_0.3rd_3_OTA_0.vd3.t13 a_21048_25880.t3 VGND.t78 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=34800,1316 d=17400,658
X51 a_3013_4521.t2 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t23 VGND.t10 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X52 a_22654_21988# 3_OTA_0.3rd_3_OTA_0.vd4.t8 a_21048_27042.t3 VGND.t78 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=34800,1316 d=17400,658
X53 VGND.t28 a_12378_15906.t32 a_12378_15906.t33 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X54 a_15996_19807# a_15996_19807# a_16084_20007# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X55 a_3013_4521.t38 a_3013_4521.t37 VGND.t47 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X56 a_3013_4521.t36 a_3013_4521.t35 VGND.t22 VGND.t21 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X57 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t27 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t9 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X58 a_6631_3101# a_6631_3101# ua[5].t3 VGND.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X59 a_3013_4521.t34 a_3013_4521.t33 VGND.t37 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X60 a_21048_27042.t11 a_21048_27042.t10 VDPWR.t41 VDPWR.t27 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=29000,1116
X61 VDPWR.t30 a_21048_25880.t8 a_21048_25880.t9 VDPWR.t29 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=29000,1116 d=14500,558
X62 a_18046_7223# ua[4].t0 VGND.t55 VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.483333 pd=3.526667 as=0 ps=0 w=3 l=5
**devattr s=34800,1316 d=34800,1316
X63 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t15 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t26 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X64 a_12378_15906.t31 a_12378_15906.t30 VGND.t23 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X65 a_16084_20007# a_15996_19807# 3_OTA_0.OTA_vref_0.vb1.t0 VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X66 3_OTA_0.3rd_3_OTA_0.vd4.t9 3_OTA_0.OTA_stage1_0.vd1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X67 ua[5].t2 a_6631_3101# a_6631_3101# VGND.t18 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X68 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t8 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t12 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X69 3_OTA_0.3rd_3_OTA_0.vd4.t2 3_OTA_0.OTA_stage1_0.vd1.t1 a_12564_25551.t2 VDPWR.t38 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X70 ua[0].t0 a_21048_27042.t12 VDPWR.t12 VDPWR.t11 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.6 l=0.35
**devattr s=30160,1156 d=30160,1156
X71 a_12378_15906.t29 a_12378_15906.t28 VGND.t31 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X72 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t1 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t11 VGND.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X73 a_15996_19807# 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t23 VDPWR.t58 VDPWR.t57 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X74 a_6719_5623# a_6631_4391# a_6719_4333# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X75 a_16084_17427# a_15996_17227# a_15996_17227# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X76 a_21048_25880.t2 3_OTA_0.3rd_3_OTA_0.vd3.t14 a_22654_21988# VGND.t77 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=34800,1316
X77 3_OTA_0.OTA_stage1_0.vd2.t1 ua[2].t1 a_3537_27009# VGND.t35 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X78 a_15996_18517# a_15996_18517# 3_OTA_0.OTA_vref_0.vb1.t5 VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X79 a_21048_27042.t2 3_OTA_0.3rd_3_OTA_0.vd4.t10 a_22654_21988# VGND.t77 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=34800,1316
X80 a_12378_15906.t41 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t13 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X81 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t13 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t25 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X82 a_16084_20007# a_15996_19807# a_15996_19807# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X83 VGND.t49 a_3013_4521.t31 a_3013_4521.t32 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X84 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t24 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t19 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X85 a_6719_6913# a_6631_6971# a_6631_6971# VGND.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X86 a_3013_4521.t30 a_3013_4521.t29 VGND.t85 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X87 a_15996_18517# 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t24 VDPWR.t56 VDPWR.t55 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X88 a_12564_25551.t10 3_OTA_0.OTA_vref_0.vb1.t7 VDPWR.t14 VDPWR.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X89 VDPWR.t69 3_OTA_0.OTA_vref_0.vb1.t8 a_12564_25551.t9 VDPWR.t68 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X90 a_21048_27042.t9 a_21048_27042.t8 VDPWR.t18 VDPWR.t17 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X91 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t7 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t23 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X92 VGND.t52 a_12378_15906.t26 a_12378_15906.t27 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X93 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t22 VDPWR.t42 VDPWR.t39 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=11600,516
X94 a_3013_4521.t47 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t22 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X95 3_OTA_0.3rd_3_OTA_0.vd3.t7 3_OTA_0.3rd_3_OTA_0.vd3.t6 VGND.t76 VGND.t69 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X96 VGND.t88 a_3013_4521.t27 a_3013_4521.t28 VGND.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X97 a_6631_5681# a_6631_5681# a_6719_5623# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X98 VGND.t14 a_12378_15906.t24 a_12378_15906.t25 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X99 VGND.t84 VGND.t83 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X100 VGND.t45 a_12378_15906.t22 a_12378_15906.t23 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X101 a_6631_3101# a_6631_3101# ua[5].t1 VGND.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X102 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t10 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t32 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X103 VGND.t12 a_3013_4521.t25 a_3013_4521.t26 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X104 VGND.t75 3_OTA_0.3rd_3_OTA_0.vd3.t4 3_OTA_0.3rd_3_OTA_0.vd3.t5 VGND.t67 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X105 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t22 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t11 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X106 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t21 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t10 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X107 a_3013_4521.t24 a_3013_4521.t23 VGND.t2 VGND.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X108 3_OTA_0.OTA_vref_0.vb a_15996_21097# a_16084_20007# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X109 a_3537_27009# ua[3].t2 3_OTA_0.OTA_stage1_0.vd1 VGND.t33 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=1.74 ps=12.58 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X110 3_OTA_0.3rd_3_OTA_0.vd4.t6 3_OTA_0.3rd_3_OTA_0.vd3.t15 VGND.t74 VGND.t73 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X111 a_15996_17227# a_15996_17227# a_16084_17427# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X112 a_3013_4521.t22 a_3013_4521.t21 VGND.t32 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X113 3_OTA_0.3rd_3_OTA_0.vd4.t1 3_OTA_0.OTA_stage1_0.vd1.t2 a_12564_25551.t3 VDPWR.t10 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X114 3_OTA_0.OTA_vref_0.vb1.t4 a_15996_18517# a_15996_18517# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X115 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t12 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 a_12378_15906.t5 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X116 a_22654_21988# 3_OTA_0.OTA_vref_0.vb VGND.t59 VGND.t58 sky130_fd_pr__nfet_01v8 ad=1.048143 pd=7.775429 as=0 ps=0 w=5.5 l=1.5
**devattr s=31900,1158 d=63800,2316
X117 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t11 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 a_12378_15906.t7 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X118 VGND.t61 a_12378_15906.t20 a_12378_15906.t21 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X119 a_6719_5623# a_6631_5681# a_6631_5681# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X120 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t9 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t2 VGND.t24 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X121 VDPWR.t54 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t25 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 VDPWR.t53 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X122 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t17 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t20 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X123 a_6631_6971# a_6631_6971# a_6719_6913# VGND.t27 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X124 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t9 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t8 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X125 a_12378_15906.t19 a_12378_15906.t18 VGND.t20 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X126 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t7 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t30 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X127 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t11 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t6 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X128 VDPWR.t33 a_18163_10306.t0 ua[1].t0 VDPWR.t31 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X129 a_21048_27042.t1 3_OTA_0.3rd_3_OTA_0.vd4.t11 a_22654_21988# VGND.t17 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=17400,658
X130 a_22654_21988# 3_OTA_0.3rd_3_OTA_0.vd4.t12 a_21048_27042.t0 VGND.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=17400,658 d=17400,658
X131 a_16084_20007# a_15996_19807# a_15996_19807# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X132 a_3537_27009# ua[2].t2 3_OTA_0.OTA_stage1_0.vd2.t0 VGND.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X133 ua[0].t2 a_25461_23684# VGND.t66 VGND.t65 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X134 VDPWR.t46 a_21048_27042.t6 a_21048_27042.t7 VDPWR.t29 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=29000,1116 d=14500,558
X135 a_15996_21097# a_15996_21097# 3_OTA_0.OTA_vref_0.vb VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=5800,258 d=5800,258
X136 a_21048_25880.t1 3_OTA_0.3rd_3_OTA_0.vd3.t16 a_22654_21988# VGND.t17 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=17400,658
X137 a_22654_21988# 3_OTA_0.3rd_3_OTA_0.vd3.t17 a_21048_25880.t0 VGND.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=17400,658 d=17400,658
X138 a_12378_15906.t3 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t10 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X139 a_16084_17427# a_15996_17227# 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t0 VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X140 a_12564_25551.t4 3_OTA_0.OTA_stage1_0.vd1.t3 3_OTA_0.3rd_3_OTA_0.vd4.t0 VDPWR.t43 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X141 VGND.t42 a_3013_4521.t19 a_3013_4521.t20 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X142 3_OTA_0.3rd_3_OTA_0.vd3.t2 3_OTA_0.OTA_stage1_0.vd2.t5 a_12564_25551.t6 VDPWR.t10 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X143 VDPWR.t26 3_OTA_0.OTA_vref_0.vb1.t9 a_12564_25551.t8 VDPWR.t25 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=81200,2916 d=40600,1458
X144 VGND.t72 3_OTA_0.3rd_3_OTA_0.vd3.t10 3_OTA_0.3rd_3_OTA_0.vd3.t11 VGND.t71 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X145 a_12378_15906.t17 a_12378_15906.t16 VGND.t25 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X146 a_12378_15906.t45 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t9 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X147 VDPWR.t21 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd2.t2 VDPWR.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X148 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t8 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 a_12378_15906.t6 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X149 a_15996_21097# 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t26 VDPWR.t52 VDPWR.t51 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X150 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t5 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t6 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X151 VGND.t29 a_12378_15906.t14 a_12378_15906.t15 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X152 a_6719_6913# a_6631_5681# a_6719_5623# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X153 3_OTA_0.OTA_vref_0.vb1.t3 a_15996_18517# a_15996_18517# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X154 VGND.t9 a_12378_15906.t12 a_12378_15906.t13 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X155 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t21 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 a_3013_4521.t9 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X156 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t4 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t3 VGND.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X157 a_21048_25880.t7 a_21048_25880.t6 VDPWR.t67 VDPWR.t17 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X158 a_6719_4333# a_6631_4391# a_6631_4391# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X159 3_OTA_0.OTA_vref_0.vb a_15996_21097# a_15996_21097# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X160 VDPWR.t65 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t23 ua[5].t5 VDPWR.t64 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X161 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t7 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 a_12378_15906.t1 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X162 a_3013_4521.t4 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t20 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X163 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t12 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t19 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X164 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t3 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t4 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X165 VGND.t51 a_3013_4521.t17 a_3013_4521.t18 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X166 a_12378_15906.t11 a_12378_15906.t10 VGND.t15 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X167 a_15996_19807# a_15996_19807# a_16084_20007# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X168 VDPWR.t20 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd1 VDPWR.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.522 ps=4.18 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X169 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t6 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 a_12378_15906.t44 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X170 VDPWR.t66 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t18 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t19 VDPWR.t15 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=5800,316 d=2900,158
X171 a_3013_4521.t45 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t19 VGND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X172 a_25461_23684# a_25461_23684# VGND.t64 VGND.t63 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X173 a_15996_17227# a_15996_17227# a_16084_17427# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X174 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t17 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t16 VDPWR.t16 VDPWR.t15 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=2900,158 d=5800,316
X175 a_3537_27009# 3_OTA_0.OTA_vref_0.vb VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.483333 pd=3.526667 as=0 ps=0 w=3 l=5
**devattr s=34800,1316 d=34800,1316
X176 a_6631_6971# a_6631_6971# a_6719_6913# VGND.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X177 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t2 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t31 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X178 VDPWR.t50 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t2 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t3 VDPWR.t48 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=5800,316 d=2900,158
X179 a_12378_15906.t46 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t5 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X180 a_6631_4391# a_6631_4391# a_6719_4333# VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X181 VDPWR.t40 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t24 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 VDPWR.t39 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X182 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t0 VDPWR.t49 VDPWR.t48 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=2900,158 d=5800,316
X183 a_12564_25551.t1 3_OTA_0.OTA_stage1_0.vd2.t6 3_OTA_0.3rd_3_OTA_0.vd3.t1 VDPWR.t43 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X184 a_3013_4521.t0 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t18 VGND.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X185 a_12378_15906.t40 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t4 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X186 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t4 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t18 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X187 a_18046_7223# ua[3].t3 ua[1].t2 VGND.t43 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X188 VDPWR.t3 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t25 a_6631_5681# VDPWR.t2 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X189 VGND.t50 a_3013_4521.t15 a_3013_4521.t16 VGND.t24 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X190 a_15996_18517# a_15996_18517# 3_OTA_0.OTA_vref_0.vb1.t2 VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X191 VDPWR.t70 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t26 a_6631_3101# VDPWR.t64 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X192 ua[5].t0 a_6631_3101# a_6631_3101# VGND.t18 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X193 a_3013_4521.t8 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t17 VGND.t19 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X194 VGND.t41 a_3013_4521.t13 a_3013_4521.t14 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X195 a_12378_15906.t9 a_12378_15906.t8 VGND.t87 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X196 a_6631_4391# a_6631_4391# a_6719_4333# VGND.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X197 VDPWR.t47 a_21048_27042.t4 a_21048_27042.t5 VDPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X198 a_25461_23684# a_21048_25880.t12 VDPWR.t5 VDPWR.t4 sky130_fd_pr__pfet_01v8_lvt ad=0.754 pd=5.78 as=0 ps=0 w=2.6 l=0.35
**devattr s=30160,1156 d=30160,1156
X199 a_12378_15906.t42 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t3 VGND.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X200 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t2 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 a_12378_15906.t2 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X201 VDPWR.t32 a_18163_10306.t0 a_18163_10306.t2 VDPWR.t31 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X202 a_12564_25551.t7 3_OTA_0.OTA_stage1_0.vd2.t7 3_OTA_0.3rd_3_OTA_0.vd3.t3 VDPWR.t37 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X203 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t16 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 a_3013_4521.t3 VGND.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X204 a_6719_6913# a_6631_6971# a_6631_6971# VGND.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X205 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t15 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 a_3013_4521.t1 VGND.t10 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X206 3_OTA_0.3rd_3_OTA_0.vd4.t5 3_OTA_0.3rd_3_OTA_0.vd3.t18 VGND.t70 VGND.t69 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X207 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t1 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t7 VGND.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X208 VGND.t82 VGND.t81 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X209 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t17 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t8 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X210 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t1 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 a_12378_15906.t4 VGND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X211 a_18046_7223# ua[2].t3 a_18163_10306.t3 VGND.t34 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X212 3_OTA_0.OTA_vref_0.vb a_15996_21097# a_15996_21097# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=11600,516
X213 3_OTA_0.OTA_vref_0.vb1.t1 a_15996_18517# a_16084_17427# VGND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X214 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t13 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t0 VGND.t89 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X215 a_21048_25880.t5 a_21048_25880.t4 VDPWR.t28 VDPWR.t27 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=29000,1116
X216 VGND.t68 3_OTA_0.3rd_3_OTA_0.vd3.t19 3_OTA_0.3rd_3_OTA_0.vd4.t4 VGND.t67 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X217 a_6719_4333# a_6631_3101# ua[5].t4 VGND.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X218 a_3013_4521.t46 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t14 VGND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
R0 3_OTA_0.3rd_3_OTA_0.vd3.n0 3_OTA_0.3rd_3_OTA_0.vd3.t14 81.6812
R1 3_OTA_0.3rd_3_OTA_0.vd3.n0 3_OTA_0.3rd_3_OTA_0.vd3.t16 81.6574
R2 3_OTA_0.3rd_3_OTA_0.vd3.n0 3_OTA_0.3rd_3_OTA_0.vd3.t17 81.6574
R3 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.3rd_3_OTA_0.vd3.t13 81.4437
R4 3_OTA_0.3rd_3_OTA_0.vd3.n2 3_OTA_0.3rd_3_OTA_0.vd3.t7 60.3532
R5 3_OTA_0.3rd_3_OTA_0.vd3.n1 3_OTA_0.3rd_3_OTA_0.vd3.t5 60.3532
R6 3_OTA_0.3rd_3_OTA_0.vd3.n3 3_OTA_0.3rd_3_OTA_0.vd3.n10 48.5755
R7 3_OTA_0.3rd_3_OTA_0.vd3.n5 3_OTA_0.3rd_3_OTA_0.vd3.t3 19.1315
R8 3_OTA_0.3rd_3_OTA_0.vd3.n5 3_OTA_0.3rd_3_OTA_0.vd3.t0 18.308
R9 3_OTA_0.3rd_3_OTA_0.vd3.n5 3_OTA_0.3rd_3_OTA_0.vd3.n6 16.2734
R10 3_OTA_0.3rd_3_OTA_0.vd3.n13 3_OTA_0.3rd_3_OTA_0.vd3.n1 14.6534
R11 3_OTA_0.3rd_3_OTA_0.vd3.n10 3_OTA_0.3rd_3_OTA_0.vd3.t11 11.6005
R12 3_OTA_0.3rd_3_OTA_0.vd3.n10 3_OTA_0.3rd_3_OTA_0.vd3.t9 11.6005
R13 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.3rd_3_OTA_0.vd3.n1 11.2227
R14 3_OTA_0.3rd_3_OTA_0.vd3.n3 3_OTA_0.3rd_3_OTA_0.vd3.n7 8.08817
R15 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.3rd_3_OTA_0.vd3.n2 7.9105
R16 3_OTA_0.3rd_3_OTA_0.vd3.n8 3_OTA_0.3rd_3_OTA_0.vd3.t6 3.58326
R17 3_OTA_0.3rd_3_OTA_0.vd3.n9 3_OTA_0.3rd_3_OTA_0.vd3.t12 3.58326
R18 3_OTA_0.3rd_3_OTA_0.vd3.n11 3_OTA_0.3rd_3_OTA_0.vd3.t15 3.58326
R19 3_OTA_0.3rd_3_OTA_0.vd3.n12 3_OTA_0.3rd_3_OTA_0.vd3.t4 3.58326
R20 3_OTA_0.3rd_3_OTA_0.vd3.n8 3_OTA_0.3rd_3_OTA_0.vd3.t18 3.58267
R21 3_OTA_0.3rd_3_OTA_0.vd3.n9 3_OTA_0.3rd_3_OTA_0.vd3.t10 3.58267
R22 3_OTA_0.3rd_3_OTA_0.vd3.n11 3_OTA_0.3rd_3_OTA_0.vd3.t8 3.58267
R23 3_OTA_0.3rd_3_OTA_0.vd3.n12 3_OTA_0.3rd_3_OTA_0.vd3.t19 3.58267
R24 3_OTA_0.3rd_3_OTA_0.vd3.n4 3_OTA_0.3rd_3_OTA_0.vd3.n13 3.54985
R25 3_OTA_0.3rd_3_OTA_0.vd3.n7 3_OTA_0.3rd_3_OTA_0.vd3.n5 2.67636
R26 3_OTA_0.3rd_3_OTA_0.vd3.n1 3_OTA_0.3rd_3_OTA_0.vd3.n12 2.60735
R27 3_OTA_0.3rd_3_OTA_0.vd3.n2 3_OTA_0.3rd_3_OTA_0.vd3.n8 2.58162
R28 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.3rd_3_OTA_0.vd3.n0 2.5555
R29 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.3rd_3_OTA_0.vd3.n7 2.29713
R30 3_OTA_0.3rd_3_OTA_0.vd3.n6 3_OTA_0.3rd_3_OTA_0.vd3.t1 1.90483
R31 3_OTA_0.3rd_3_OTA_0.vd3.n6 3_OTA_0.3rd_3_OTA_0.vd3.t2 1.90483
R32 3_OTA_0.3rd_3_OTA_0.vd3.n2 3_OTA_0.3rd_3_OTA_0.vd3.n4 1.69798
R33 3_OTA_0.3rd_3_OTA_0.vd3.n13 3_OTA_0.3rd_3_OTA_0.vd3.n11 1.61224
R34 3_OTA_0.3rd_3_OTA_0.vd3.n4 3_OTA_0.3rd_3_OTA_0.vd3.n9 1.61224
R35 3_OTA_0.3rd_3_OTA_0.vd3.n4 3_OTA_0.3rd_3_OTA_0.vd3.n3 1.22519
R36 VGND.n743 VGND.n249 5.69811e+06
R37 VGND.n532 VGND.n531 2.37903e+06
R38 VGND.n298 VGND.n249 1.38761e+06
R39 VGND.n531 VGND.n530 882739
R40 VGND.n514 VGND.n509 702439
R41 VGND.n526 VGND.n509 498262
R42 VGND.n527 VGND.n526 496062
R43 VGND.n530 VGND.n529 434133
R44 VGND.n528 VGND.n527 349800
R45 VGND.n360 VGND.n335 156933
R46 VGND.n441 VGND.n335 128213
R47 VGND.n529 VGND.n528 123200
R48 VGND.n525 VGND.n524 45325.3
R49 VGND.n763 VGND.n762 38916.1
R50 VGND.n409 VGND.n385 27614.8
R51 VGND.n453 VGND.n385 27609
R52 VGND.n409 VGND.n386 27609
R53 VGND.n453 VGND.n386 27603.2
R54 VGND.n794 VGND.n7 26954.2
R55 VGND.n794 VGND.n6 26954.2
R56 VGND.n745 VGND.n234 26954.2
R57 VGND.n757 VGND.n234 26954.2
R58 VGND.n796 VGND.n6 26948.4
R59 VGND.n796 VGND.n7 26948.4
R60 VGND.n745 VGND.n236 26948.4
R61 VGND.n757 VGND.n236 26948.4
R62 VGND.n436 VGND.n388 25442
R63 VGND.n436 VGND.n389 25442
R64 VGND.n309 VGND.n305 25442
R65 VGND.n496 VGND.n309 25442
R66 VGND.n448 VGND.n388 25436.2
R67 VGND.n448 VGND.n389 25436.2
R68 VGND.n497 VGND.n305 25436.2
R69 VGND.n497 VGND.n496 25436.2
R70 VGND.n529 VGND.n297 24244.5
R71 VGND.n441 VGND.n440 24216.7
R72 VGND.n760 VGND.t8 21212.8
R73 VGND.n528 VGND.n298 20643.3
R74 VGND.n742 VGND.n250 17753.2
R75 VGND.n742 VGND.n251 17753.2
R76 VGND.n738 VGND.n250 17753.2
R77 VGND.n738 VGND.n251 17753.2
R78 VGND.n523 VGND.n512 17753.2
R79 VGND.n523 VGND.n515 17753.2
R80 VGND.n518 VGND.n512 17753.2
R81 VGND.n518 VGND.n515 17753.2
R82 VGND.n442 VGND.n437 16119.1
R83 VGND.n761 VGND.t5 15479.6
R84 VGND.n517 VGND.t1 13323.7
R85 VGND.n356 VGND.n336 12277.7
R86 VGND.n468 VGND.n336 12277.7
R87 VGND.n356 VGND.n338 12277.7
R88 VGND.n468 VGND.n338 12277.7
R89 VGND.n360 VGND.n310 11383.3
R90 VGND.n528 VGND.n508 10329.2
R91 VGND.n451 VGND.t8 10154.9
R92 VGND.n762 VGND.n761 8959.58
R93 VGND.n531 VGND.n232 8257.79
R94 VGND.n443 VGND.n442 7054.95
R95 VGND.n353 VGND.n333 6732.77
R96 VGND.n471 VGND.n333 6732.77
R97 VGND.n353 VGND.n334 6732.77
R98 VGND.n471 VGND.n334 6732.77
R99 VGND.n445 VGND.n392 6275.03
R100 VGND.n393 VGND.n392 6275.03
R101 VGND.n445 VGND.n444 6275.03
R102 VGND.n444 VGND.n393 6275.03
R103 VGND.n500 VGND.n299 6275.03
R104 VGND.n507 VGND.n299 6275.03
R105 VGND.n500 VGND.n300 6275.03
R106 VGND.n507 VGND.n300 6275.03
R107 VGND.t18 VGND.t21 5886.96
R108 VGND.n452 VGND.n451 5653.83
R109 VGND.t5 VGND.n230 5382.74
R110 VGND.n491 VGND.n312 4519.41
R111 VGND.n491 VGND.n313 4519.41
R112 VGND.n358 VGND.n312 4519.41
R113 VGND.n358 VGND.n313 4519.41
R114 VGND.t3 VGND.t16 4306.23
R115 VGND.n760 VGND.n759 4090.89
R116 VGND.n451 VGND.n450 4053.37
R117 VGND.t3 VGND.n245 4004.26
R118 VGND.t5 VGND.n51 4004.26
R119 VGND.n761 VGND.n760 3745.57
R120 VGND.n235 VGND.n231 3636.37
R121 VGND.n364 VGND.n343 3412.74
R122 VGND.n366 VGND.n343 3412.74
R123 VGND.n364 VGND.n344 3406.94
R124 VGND.n366 VGND.n344 3406.94
R125 VGND.n532 VGND.n249 3402.79
R126 VGND.t73 VGND.t67 3214.17
R127 VGND.n94 VGND.n93 3100.52
R128 VGND.n225 VGND.n8 3064.3
R129 VGND.n494 VGND.n493 3057.55
R130 VGND.n441 VGND.n310 3019.08
R131 VGND.n524 VGND.t39 2995.18
R132 VGND.n517 VGND.t39 2906.83
R133 VGND.t1 VGND.n511 2812.74
R134 VGND.n513 VGND.t21 2381.06
R135 VGND.n93 VGND.n64 2051.81
R136 VGND.n155 VGND.n64 2051.81
R137 VGND.n156 VGND.n155 2051.81
R138 VGND.n158 VGND.n156 2051.81
R139 VGND.n158 VGND.n157 2051.81
R140 VGND.n172 VGND.n171 2051.81
R141 VGND.n173 VGND.n172 2051.81
R142 VGND.n173 VGND.n56 2051.81
R143 VGND.n182 VGND.n56 2051.81
R144 VGND.n183 VGND.n182 2051.81
R145 VGND.n763 VGND.n183 2051.81
R146 VGND.n452 VGND.t67 1975.27
R147 VGND.n442 VGND.n441 1964.94
R148 VGND.n488 VGND.n487 1960.4
R149 VGND.n758 VGND.n233 1584.56
R150 VGND.n437 VGND.t30 1579.6
R151 VGND.n450 VGND.n449 1546.15
R152 VGND.n439 VGND.t71 1508.37
R153 VGND.n157 VGND.t84 1390.67
R154 VGND.t35 VGND.n395 1326.04
R155 VGND.n395 VGND.t62 1324.96
R156 VGND.n766 VGND.n53 1305.6
R157 VGND.n699 VGND.n698 1305.6
R158 VGND.n440 VGND.t73 1287
R159 VGND.n741 VGND.n244 1245.36
R160 VGND.n514 VGND.n513 1243.41
R161 VGND.n759 VGND.n758 1221.6
R162 VGND.n116 VGND.n95 1168.03
R163 VGND.n525 VGND.t6 1166.51
R164 VGND.n514 VGND.t89 1121.63
R165 VGND.n493 VGND.n310 1115.47
R166 VGND.n759 VGND.n232 1100
R167 VGND.n493 VGND.n492 914.144
R168 VGND.n455 VGND.n383 903.91
R169 VGND.t48 VGND.n494 675.149
R170 VGND.n498 VGND.t43 675.149
R171 VGND.n745 VGND.n744 661.352
R172 VGND.n171 VGND.t84 661.14
R173 VGND.n235 VGND.t8 651.01
R174 VGND.t3 VGND.n246 647.059
R175 VGND.n760 VGND.n231 637.181
R176 VGND.n737 VGND.n736 635.574
R177 VGND.n119 VGND.n86 588.759
R178 VGND.n90 VGND.n89 588.759
R179 VGND.n676 VGND.n675 588.759
R180 VGND.n560 VGND.n538 588.759
R181 VGND.n355 VGND.n339 588.515
R182 VGND.n95 VGND.n86 585
R183 VGND.n224 VGND.n223 585
R184 VGND.n223 VGND.n222 585
R185 VGND.n23 VGND.n20 585
R186 VGND.n20 VGND.n19 585
R187 VGND.n778 VGND.n777 585
R188 VGND.n779 VGND.n778 585
R189 VGND.n21 VGND.n18 585
R190 VGND.n780 VGND.n18 585
R191 VGND.n783 VGND.n782 585
R192 VGND.n782 VGND.n781 585
R193 VGND.n103 VGND.n17 585
R194 VGND.n99 VGND.n17 585
R195 VGND.n102 VGND.n101 585
R196 VGND.n101 VGND.n100 585
R197 VGND.n108 VGND.n97 585
R198 VGND.n97 VGND.n96 585
R199 VGND.n113 VGND.n112 585
R200 VGND.n114 VGND.n113 585
R201 VGND.n88 VGND.n87 585
R202 VGND.n115 VGND.n88 585
R203 VGND.n118 VGND.n117 585
R204 VGND.n117 VGND.n116 585
R205 VGND.n69 VGND.n67 585
R206 VGND.n144 VGND.n143 585
R207 VGND.n77 VGND.n70 585
R208 VGND.n139 VGND.n138 585
R209 VGND.n82 VGND.n76 585
R210 VGND.n133 VGND.n132 585
R211 VGND.n125 VGND.n83 585
R212 VGND.n127 VGND.n126 585
R213 VGND.n85 VGND.n84 585
R214 VGND.n120 VGND.n73 585
R215 VGND.n141 VGND.n73 585
R216 VGND.n181 VGND.n180 585
R217 VGND.n182 VGND.n181 585
R218 VGND.n178 VGND.n57 585
R219 VGND.n57 VGND.n56 585
R220 VGND.n175 VGND.n174 585
R221 VGND.n174 VGND.n173 585
R222 VGND.n166 VGND.n59 585
R223 VGND.n172 VGND.n59 585
R224 VGND.n170 VGND.n169 585
R225 VGND.n171 VGND.n170 585
R226 VGND.n61 VGND.n60 585
R227 VGND.n157 VGND.n60 585
R228 VGND.n160 VGND.n159 585
R229 VGND.n159 VGND.n158 585
R230 VGND.n149 VGND.n63 585
R231 VGND.n156 VGND.n63 585
R232 VGND.n154 VGND.n153 585
R233 VGND.n155 VGND.n154 585
R234 VGND.n66 VGND.n65 585
R235 VGND.n65 VGND.n64 585
R236 VGND.n92 VGND.n91 585
R237 VGND.n93 VGND.n92 585
R238 VGND.n765 VGND.n764 585
R239 VGND.n764 VGND.n763 585
R240 VGND.n55 VGND.n54 585
R241 VGND.n183 VGND.n55 585
R242 VGND.n52 VGND.n51 585
R243 VGND.n228 VGND.n227 585
R244 VGND.n228 VGND.n51 585
R245 VGND.n219 VGND.n186 585
R246 VGND.n216 VGND.n215 585
R247 VGND.n213 VGND.n188 585
R248 VGND.n211 VGND.n210 585
R249 VGND.n202 VGND.n189 585
R250 VGND.n201 VGND.n200 585
R251 VGND.n198 VGND.n196 585
R252 VGND.n191 VGND.n50 585
R253 VGND.n771 VGND.n770 585
R254 VGND.n230 VGND.n229 585
R255 VGND.n221 VGND.n184 585
R256 VGND.n702 VGND.n245 585
R257 VGND.n701 VGND.n700 585
R258 VGND.n701 VGND.n233 585
R259 VGND.n281 VGND.n280 585
R260 VGND.n694 VGND.n280 585
R261 VGND.n706 VGND.n705 585
R262 VGND.n278 VGND.n275 585
R263 VGND.n272 VGND.n270 585
R264 VGND.n714 VGND.n713 585
R265 VGND.n717 VGND.n716 585
R266 VGND.n269 VGND.n266 585
R267 VGND.n262 VGND.n260 585
R268 VGND.n725 VGND.n724 585
R269 VGND.n727 VGND.n259 585
R270 VGND.n728 VGND.n254 585
R271 VGND.n728 VGND.n245 585
R272 VGND.n697 VGND.n696 585
R273 VGND.n696 VGND.n695 585
R274 VGND.n287 VGND.n283 585
R275 VGND.n693 VGND.n283 585
R276 VGND.n691 VGND.n690 585
R277 VGND.n692 VGND.n691 585
R278 VGND.n290 VGND.n285 585
R279 VGND.n285 VGND.n284 585
R280 VGND.n681 VGND.n680 585
R281 VGND.n680 VGND.n679 585
R282 VGND.n294 VGND.n293 585
R283 VGND.n295 VGND.n294 585
R284 VGND.n637 VGND.n636 585
R285 VGND.n638 VGND.n637 585
R286 VGND.n565 VGND.n559 585
R287 VGND.n639 VGND.n559 585
R288 VGND.n642 VGND.n641 585
R289 VGND.n641 VGND.n640 585
R290 VGND.n558 VGND.n556 585
R291 VGND.n564 VGND.n558 585
R292 VGND.n562 VGND.n561 585
R293 VGND.n563 VGND.n562 585
R294 VGND.n674 VGND.n540 585
R295 VGND.n543 VGND.n539 585
R296 VGND.n678 VGND.n539 585
R297 VGND.n669 VGND.n668 585
R298 VGND.n661 VGND.n546 585
R299 VGND.n663 VGND.n662 585
R300 VGND.n654 VGND.n548 585
R301 VGND.n656 VGND.n655 585
R302 VGND.n647 VGND.n551 585
R303 VGND.n649 VGND.n648 585
R304 VGND.n554 VGND.n553 585
R305 VGND.n678 VGND.n538 585
R306 VGND.n730 VGND.n729 585
R307 VGND.n731 VGND.n257 585
R308 VGND.n734 VGND.n733 585
R309 VGND.n733 VGND.n732 585
R310 VGND.n591 VGND.n256 585
R311 VGND.n258 VGND.n256 585
R312 VGND.n626 VGND.n625 585
R313 VGND.n627 VGND.n626 585
R314 VGND.n589 VGND.n587 585
R315 VGND.n628 VGND.n587 585
R316 VGND.n631 VGND.n630 585
R317 VGND.n630 VGND.n629 585
R318 VGND.n594 VGND.n586 585
R319 VGND.n610 VGND.n586 585
R320 VGND.n613 VGND.n612 585
R321 VGND.n612 VGND.n611 585
R322 VGND.n609 VGND.n597 585
R323 VGND.n609 VGND.n248 585
R324 VGND.n608 VGND.n603 585
R325 VGND.n608 VGND.n607 585
R326 VGND.n599 VGND.n598 585
R327 VGND.n606 VGND.n598 585
R328 VGND.n542 VGND.n541 585
R329 VGND.n605 VGND.n541 585
R330 VGND.n495 VGND.t13 566.775
R331 VGND.n495 VGND.t34 566.314
R332 VGND.n408 VGND.n335 562.178
R333 VGND.n377 VGND.n339 512.625
R334 VGND.n116 VGND.n115 502.538
R335 VGND.n115 VGND.n114 502.538
R336 VGND.n114 VGND.n96 502.538
R337 VGND.n100 VGND.n96 502.538
R338 VGND.n100 VGND.n99 502.538
R339 VGND.n781 VGND.n780 502.538
R340 VGND.n780 VGND.n779 502.538
R341 VGND.n779 VGND.n19 502.538
R342 VGND.n222 VGND.n19 502.538
R343 VGND.n222 VGND.n184 502.538
R344 VGND.n230 VGND.n184 502.538
R345 VGND.t56 VGND.n387 493.086
R346 VGND.t56 VGND.n443 493.086
R347 VGND.n744 VGND.t3 443.885
R348 VGND.n744 VGND.t8 440.897
R349 VGND.n449 VGND.n387 391.663
R350 VGND.n408 VGND.t69 382.955
R351 VGND.n440 VGND.n439 356.233
R352 VGND.t69 VGND.n298 341.902
R353 VGND.n99 VGND.t84 340.61
R354 VGND.t82 VGND.n678 331.916
R355 VGND.n71 VGND.t84 322.904
R356 VGND.t82 VGND.n245 319.149
R357 VGND.n51 VGND.t84 319.149
R358 VGND.n95 VGND.n94 319.084
R359 VGND.n435 VGND.n396 307.036
R360 VGND.n308 VGND.n307 307.036
R361 VGND.n730 VGND.n246 305.255
R362 VGND.n491 VGND.n490 292.5
R363 VGND.n492 VGND.n491 292.5
R364 VGND.n358 VGND.n315 292.5
R365 VGND.n359 VGND.n358 292.5
R366 VGND.n522 VGND.n521 281.336
R367 VGND.n740 VGND.n739 281.336
R368 VGND.n522 VGND.n516 281.243
R369 VGND.n741 VGND.n740 281.243
R370 VGND.n346 VGND.n318 270.709
R371 VGND.n421 VGND.n420 262.366
R372 VGND.n645 VGND.n644 258.334
R373 VGND.n147 VGND.n146 258.334
R374 VGND.n676 VGND.n541 257.466
R375 VGND.n117 VGND.n86 257.466
R376 VGND.n396 VGND.n390 256.805
R377 VGND.n307 VGND.n306 256.805
R378 VGND.n797 VGND.n5 255.26
R379 VGND.n747 VGND.n746 255.26
R380 VGND.n141 VGND.n72 254.34
R381 VGND.n142 VGND.n141 254.34
R382 VGND.n141 VGND.n140 254.34
R383 VGND.n141 VGND.n75 254.34
R384 VGND.n141 VGND.n74 254.34
R385 VGND.n768 VGND.n767 254.34
R386 VGND.n769 VGND.n51 254.34
R387 VGND.n214 VGND.n51 254.34
R388 VGND.n212 VGND.n51 254.34
R389 VGND.n199 VGND.n51 254.34
R390 VGND.n197 VGND.n51 254.34
R391 VGND.n225 VGND.n185 254.34
R392 VGND.n703 VGND.n279 254.34
R393 VGND.n704 VGND.n245 254.34
R394 VGND.n277 VGND.n245 254.34
R395 VGND.n715 VGND.n245 254.34
R396 VGND.n268 VGND.n245 254.34
R397 VGND.n726 VGND.n245 254.34
R398 VGND.n678 VGND.n677 254.34
R399 VGND.n678 VGND.n534 254.34
R400 VGND.n678 VGND.n535 254.34
R401 VGND.n678 VGND.n536 254.34
R402 VGND.n678 VGND.n537 254.34
R403 VGND.n736 VGND.n253 254.34
R404 VGND.n419 VGND.n418 252.304
R405 VGND.n562 VGND.n538 249.663
R406 VGND.n92 VGND.n89 249.663
R407 VGND.t71 VGND.n298 240.571
R408 VGND.n410 VGND.n381 223.468
R409 VGND.n773 VGND.n45 221.667
R410 VGND.n429 VGND.n428 216.017
R411 VGND.n506 VGND.n301 216.017
R412 VGND.n94 VGND.n71 215.269
R413 VGND.n499 VGND.t54 210.755
R414 VGND.n508 VGND.t54 210.755
R415 VGND.n678 VGND.n533 208.512
R416 VGND.n48 VGND.n47 200.388
R417 VGND.n756 VGND.n237 200.388
R418 VGND.n220 VGND.n25 185
R419 VGND.n776 VGND.n775 185
R420 VGND.n24 VGND.n22 185
R421 VGND.n37 VGND.n16 185
R422 VGND.n36 VGND.n15 185
R423 VGND.n105 VGND.n104 185
R424 VGND.n107 VGND.n106 185
R425 VGND.n111 VGND.n110 185
R426 VGND.n109 VGND.n98 185
R427 VGND.n146 VGND.n145 185
R428 VGND.n78 VGND.n68 185
R429 VGND.n80 VGND.n79 185
R430 VGND.n137 VGND.n136 185
R431 VGND.n135 VGND.n134 185
R432 VGND.n131 VGND.n130 185
R433 VGND.n129 VGND.n128 185
R434 VGND.n124 VGND.n123 185
R435 VGND.n122 VGND.n121 185
R436 VGND.n179 VGND.n45 185
R437 VGND.n177 VGND.n176 185
R438 VGND.n58 VGND.n39 185
R439 VGND.t83 VGND.n39 185
R440 VGND.n168 VGND.n167 185
R441 VGND.n165 VGND.n164 185
R442 VGND.n163 VGND.n162 185
R443 VGND.n150 VGND.n62 185
R444 VGND.n152 VGND.n151 185
R445 VGND.n148 VGND.n147 185
R446 VGND.n218 VGND.n217 185
R447 VGND.n207 VGND.n187 185
R448 VGND.n209 VGND.n208 185
R449 VGND.n206 VGND.n205 185
R450 VGND.n204 VGND.n203 185
R451 VGND.n193 VGND.n190 185
R452 VGND.n195 VGND.n194 185
R453 VGND.n49 VGND.n46 185
R454 VGND.n773 VGND.n772 185
R455 VGND.t83 VGND.n773 185
R456 VGND.n276 VGND.n274 185
R457 VGND.n708 VGND.n707 185
R458 VGND.n710 VGND.n273 185
R459 VGND.n712 VGND.n711 185
R460 VGND.n267 VGND.n265 185
R461 VGND.n719 VGND.n718 185
R462 VGND.n721 VGND.n264 185
R463 VGND.n723 VGND.n722 185
R464 VGND.n592 VGND.n261 185
R465 VGND.n593 VGND.n255 185
R466 VGND.n593 VGND.t81 185
R467 VGND.n624 VGND.n623 185
R468 VGND.n621 VGND.n590 185
R469 VGND.n620 VGND.n585 185
R470 VGND.n618 VGND.n584 185
R471 VGND.n617 VGND.n595 185
R472 VGND.n615 VGND.n614 185
R473 VGND.n602 VGND.n596 185
R474 VGND.n596 VGND.t81 185
R475 VGND.n601 VGND.n600 185
R476 VGND.n673 VGND.n672 185
R477 VGND.n671 VGND.n670 185
R478 VGND.n667 VGND.n666 185
R479 VGND.n665 VGND.n664 185
R480 VGND.n660 VGND.n659 185
R481 VGND.n658 VGND.n657 185
R482 VGND.n653 VGND.n652 185
R483 VGND.n651 VGND.n650 185
R484 VGND.n646 VGND.n645 185
R485 VGND.n289 VGND.n282 185
R486 VGND.n689 VGND.n688 185
R487 VGND.n686 VGND.n286 185
R488 VGND.n685 VGND.n291 185
R489 VGND.n683 VGND.n682 185
R490 VGND.n570 VGND.n292 185
R491 VGND.n569 VGND.n568 185
R492 VGND.n566 VGND.n557 185
R493 VGND.n644 VGND.n643 185
R494 VGND.n447 VGND.n390 184.031
R495 VGND.n306 VGND.n304 184.031
R496 VGND.n435 VGND.n434 177.084
R497 VGND.n308 VGND.n303 177.084
R498 VGND.n598 VGND.n541 175.546
R499 VGND.n608 VGND.n598 175.546
R500 VGND.n609 VGND.n608 175.546
R501 VGND.n612 VGND.n609 175.546
R502 VGND.n612 VGND.n586 175.546
R503 VGND.n630 VGND.n586 175.546
R504 VGND.n630 VGND.n587 175.546
R505 VGND.n626 VGND.n587 175.546
R506 VGND.n626 VGND.n256 175.546
R507 VGND.n733 VGND.n256 175.546
R508 VGND.n733 VGND.n257 175.546
R509 VGND.n540 VGND.n539 175.546
R510 VGND.n668 VGND.n539 175.546
R511 VGND.n662 VGND.n661 175.546
R512 VGND.n655 VGND.n654 175.546
R513 VGND.n648 VGND.n647 175.546
R514 VGND.n553 VGND.n538 175.546
R515 VGND.n562 VGND.n558 175.546
R516 VGND.n641 VGND.n558 175.546
R517 VGND.n641 VGND.n559 175.546
R518 VGND.n637 VGND.n559 175.546
R519 VGND.n637 VGND.n294 175.546
R520 VGND.n680 VGND.n294 175.546
R521 VGND.n680 VGND.n285 175.546
R522 VGND.n691 VGND.n285 175.546
R523 VGND.n691 VGND.n283 175.546
R524 VGND.n696 VGND.n283 175.546
R525 VGND.n696 VGND.n280 175.546
R526 VGND.n701 VGND.n280 175.546
R527 VGND.n728 VGND.n727 175.546
R528 VGND.n725 VGND.n260 175.546
R529 VGND.n716 VGND.n269 175.546
R530 VGND.n714 VGND.n270 175.546
R531 VGND.n705 VGND.n278 175.546
R532 VGND.n92 VGND.n65 175.546
R533 VGND.n154 VGND.n65 175.546
R534 VGND.n154 VGND.n63 175.546
R535 VGND.n159 VGND.n63 175.546
R536 VGND.n159 VGND.n60 175.546
R537 VGND.n170 VGND.n60 175.546
R538 VGND.n170 VGND.n59 175.546
R539 VGND.n174 VGND.n59 175.546
R540 VGND.n174 VGND.n57 175.546
R541 VGND.n181 VGND.n57 175.546
R542 VGND.n181 VGND.n55 175.546
R543 VGND.n764 VGND.n55 175.546
R544 VGND.n770 VGND.n50 175.546
R545 VGND.n200 VGND.n198 175.546
R546 VGND.n211 VGND.n189 175.546
R547 VGND.n215 VGND.n213 175.546
R548 VGND.n228 VGND.n186 175.546
R549 VGND.n117 VGND.n88 175.546
R550 VGND.n113 VGND.n88 175.546
R551 VGND.n113 VGND.n97 175.546
R552 VGND.n101 VGND.n97 175.546
R553 VGND.n101 VGND.n17 175.546
R554 VGND.n782 VGND.n17 175.546
R555 VGND.n782 VGND.n18 175.546
R556 VGND.n778 VGND.n18 175.546
R557 VGND.n778 VGND.n20 175.546
R558 VGND.n223 VGND.n20 175.546
R559 VGND.n223 VGND.n221 175.546
R560 VGND.n143 VGND.n69 175.546
R561 VGND.n139 VGND.n70 175.546
R562 VGND.n132 VGND.n76 175.546
R563 VGND.n126 VGND.n125 175.546
R564 VGND.n84 VGND.n73 175.546
R565 VGND.n86 VGND.n73 175.546
R566 VGND.n359 VGND.n357 170.339
R567 VGND.n458 VGND.n457 169.446
R568 VGND.n499 VGND.n498 167.405
R569 VGND.n593 VGND.n592 163.333
R570 VGND.n217 VGND.n25 163.333
R571 VGND.n781 VGND.t84 161.929
R572 VGND.n704 VGND.n703 152.643
R573 VGND.n769 VGND.n768 152.643
R574 VGND.n600 VGND.n596 150
R575 VGND.n615 VGND.n596 150
R576 VGND.n618 VGND.n617 150
R577 VGND.n621 VGND.n620 150
R578 VGND.n623 VGND.n593 150
R579 VGND.n672 VGND.n671 150
R580 VGND.n666 VGND.n665 150
R581 VGND.n659 VGND.n658 150
R582 VGND.n652 VGND.n651 150
R583 VGND.n568 VGND.n566 150
R584 VGND.n683 VGND.n292 150
R585 VGND.n686 VGND.n685 150
R586 VGND.n688 VGND.n289 150
R587 VGND.n722 VGND.n721 150
R588 VGND.n719 VGND.n265 150
R589 VGND.n711 VGND.n710 150
R590 VGND.n708 VGND.n274 150
R591 VGND.n79 VGND.n78 150
R592 VGND.n136 VGND.n135 150
R593 VGND.n130 VGND.n129 150
R594 VGND.n123 VGND.n122 150
R595 VGND.n151 VGND.n150 150
R596 VGND.n164 VGND.n163 150
R597 VGND.n167 VGND.n39 150
R598 VGND.n176 VGND.n39 150
R599 VGND.n773 VGND.n46 150
R600 VGND.n194 VGND.n193 150
R601 VGND.n205 VGND.n204 150
R602 VGND.n208 VGND.n207 150
R603 VGND.n110 VGND.n109 150
R604 VGND.n106 VGND.n105 150
R605 VGND.n37 VGND.n36 150
R606 VGND.n775 VGND.n24 150
R607 VGND.n490 VGND.n489 149.538
R608 VGND.n520 VGND.n5 147.642
R609 VGND.n746 VGND.n244 147.642
R610 VGND.n729 VGND.n728 146.287
R611 VGND.n229 VGND.n228 146.287
R612 VGND.n360 VGND.n359 143.072
R613 VGND.t77 VGND.t0 140.315
R614 VGND.n702 VGND.n701 138.486
R615 VGND.n764 VGND.n52 138.486
R616 VGND.n470 VGND.t17 138.477
R617 VGND.n805 VGND.n4 137.462
R618 VGND.n755 VGND.n238 137.462
R619 VGND.n605 VGND.n604 130.4
R620 VGND.n489 VGND.n488 126.4
R621 VGND.n563 VGND.n533 123.46
R622 VGND.n805 VGND.n804 122.373
R623 VGND.n748 VGND.n238 122.373
R624 VGND.n467 VGND.n466 113.549
R625 VGND.n467 VGND.n377 109.558
R626 VGND.n486 VGND.n317 104.918
R627 VGND.t78 VGND.n469 103.858
R628 VGND.n344 VGND.n342 97.5005
R629 VGND.n361 VGND.n344 97.5005
R630 VGND.n362 VGND.n343 97.5005
R631 VGND.n343 VGND.n311 97.5005
R632 VGND.n357 VGND.n354 94.667
R633 VGND.n433 VGND.n391 89.9525
R634 VGND.n503 VGND.n502 89.9525
R635 VGND.n340 VGND.t66 89.2211
R636 VGND.n340 VGND.t64 89.0687
R637 VGND.n606 VGND.n605 88.9093
R638 VGND.n607 VGND.n606 88.9093
R639 VGND.n611 VGND.n248 88.9093
R640 VGND.n611 VGND.n610 88.9093
R641 VGND.n629 VGND.n628 88.9093
R642 VGND.n628 VGND.n627 88.9093
R643 VGND.n627 VGND.n258 88.9093
R644 VGND.n732 VGND.n258 88.9093
R645 VGND.n732 VGND.n731 88.9093
R646 VGND.n731 VGND.n730 88.9093
R647 VGND.n564 VGND.n563 83.5448
R648 VGND.n640 VGND.n564 83.5448
R649 VGND.n640 VGND.n639 83.5448
R650 VGND.n639 VGND.n638 83.5448
R651 VGND.n638 VGND.n295 83.5448
R652 VGND.n679 VGND.n284 83.5448
R653 VGND.n692 VGND.n284 83.5448
R654 VGND.n693 VGND.n692 83.5448
R655 VGND.n695 VGND.n693 83.5448
R656 VGND.n695 VGND.n694 83.5448
R657 VGND.n694 VGND.n233 83.5448
R658 VGND.n515 VGND.t18 81.0238
R659 VGND.n526 VGND.n525 79.3569
R660 VGND.n729 VGND.n253 76.3222
R661 VGND.n677 VGND.n676 76.3222
R662 VGND.n668 VGND.n534 76.3222
R663 VGND.n662 VGND.n535 76.3222
R664 VGND.n655 VGND.n536 76.3222
R665 VGND.n648 VGND.n537 76.3222
R666 VGND.n726 VGND.n725 76.3222
R667 VGND.n269 VGND.n268 76.3222
R668 VGND.n715 VGND.n714 76.3222
R669 VGND.n278 VGND.n277 76.3222
R670 VGND.n703 VGND.n702 76.3222
R671 VGND.n197 VGND.n50 76.3222
R672 VGND.n200 VGND.n199 76.3222
R673 VGND.n212 VGND.n211 76.3222
R674 VGND.n215 VGND.n214 76.3222
R675 VGND.n229 VGND.n185 76.3222
R676 VGND.n72 VGND.n69 76.3222
R677 VGND.n143 VGND.n142 76.3222
R678 VGND.n140 VGND.n139 76.3222
R679 VGND.n132 VGND.n75 76.3222
R680 VGND.n126 VGND.n74 76.3222
R681 VGND.n142 VGND.n70 76.3222
R682 VGND.n140 VGND.n76 76.3222
R683 VGND.n125 VGND.n75 76.3222
R684 VGND.n84 VGND.n74 76.3222
R685 VGND.n89 VGND.n72 76.3222
R686 VGND.n768 VGND.n52 76.3222
R687 VGND.n214 VGND.n186 76.3222
R688 VGND.n213 VGND.n212 76.3222
R689 VGND.n199 VGND.n189 76.3222
R690 VGND.n198 VGND.n197 76.3222
R691 VGND.n770 VGND.n769 76.3222
R692 VGND.n221 VGND.n185 76.3222
R693 VGND.n705 VGND.n704 76.3222
R694 VGND.n277 VGND.n270 76.3222
R695 VGND.n716 VGND.n715 76.3222
R696 VGND.n268 VGND.n260 76.3222
R697 VGND.n727 VGND.n726 76.3222
R698 VGND.n677 VGND.n540 76.3222
R699 VGND.n661 VGND.n534 76.3222
R700 VGND.n654 VGND.n535 76.3222
R701 VGND.n647 VGND.n536 76.3222
R702 VGND.n553 VGND.n537 76.3222
R703 VGND.n257 VGND.n253 76.3222
R704 VGND.n672 VGND.n544 74.5978
R705 VGND.n122 VGND.n32 74.5978
R706 VGND.n109 VGND.n32 74.5978
R707 VGND.n600 VGND.n544 74.5978
R708 VGND.n363 VGND.n362 73.0981
R709 VGND.n345 VGND.t17 72.6088
R710 VGND.n289 VGND.n288 69.3109
R711 VGND.n288 VGND.n274 69.3109
R712 VGND.n418 VGND.n410 69.0601
R713 VGND.n521 VGND.n520 68.6416
R714 VGND.n774 VGND.t83 65.8183
R715 VGND.t83 VGND.n38 65.8183
R716 VGND.t83 VGND.n34 65.8183
R717 VGND.t83 VGND.n27 65.8183
R718 VGND.t83 VGND.n28 65.8183
R719 VGND.t83 VGND.n29 65.8183
R720 VGND.t83 VGND.n30 65.8183
R721 VGND.t83 VGND.n31 65.8183
R722 VGND.t83 VGND.n40 65.8183
R723 VGND.t83 VGND.n35 65.8183
R724 VGND.t83 VGND.n33 65.8183
R725 VGND.t83 VGND.n26 65.8183
R726 VGND.t83 VGND.n41 65.8183
R727 VGND.t83 VGND.n42 65.8183
R728 VGND.t83 VGND.n43 65.8183
R729 VGND.t83 VGND.n44 65.8183
R730 VGND.n709 VGND.t81 65.8183
R731 VGND.n271 VGND.t81 65.8183
R732 VGND.n720 VGND.t81 65.8183
R733 VGND.t81 VGND.n263 65.8183
R734 VGND.n622 VGND.t81 65.8183
R735 VGND.n619 VGND.t81 65.8183
R736 VGND.n616 VGND.t81 65.8183
R737 VGND.n545 VGND.t81 65.8183
R738 VGND.n547 VGND.t81 65.8183
R739 VGND.n549 VGND.t81 65.8183
R740 VGND.n552 VGND.t81 65.8183
R741 VGND.n687 VGND.t81 65.8183
R742 VGND.n684 VGND.t81 65.8183
R743 VGND.n567 VGND.t81 65.8183
R744 VGND.n555 VGND.t81 65.8183
R745 VGND.n521 VGND.n515 65.0005
R746 VGND.n516 VGND.n512 65.0005
R747 VGND.n512 VGND.n296 65.0005
R748 VGND.n367 VGND.n366 65.0005
R749 VGND.n366 VGND.n365 65.0005
R750 VGND.n364 VGND.n363 65.0005
R751 VGND.n365 VGND.n364 65.0005
R752 VGND.n739 VGND.n738 65.0005
R753 VGND.n738 VGND.n247 65.0005
R754 VGND.n742 VGND.n741 65.0005
R755 VGND.n743 VGND.n742 65.0005
R756 VGND.t16 VGND.n248 62.2367
R757 VGND.t0 VGND.t58 62.1924
R758 VGND.n610 VGND.t82 60.2609
R759 VGND.n365 VGND.t65 59.9007
R760 VGND.n365 VGND.t63 58.5695
R761 VGND.n288 VGND.t81 57.8461
R762 VGND.t82 VGND.n295 56.625
R763 VGND.n363 VGND.n342 56.241
R764 VGND.t83 VGND.n32 55.2026
R765 VGND.n544 VGND.t81 55.2026
R766 VGND.t65 VGND.n311 54.2434
R767 VGND.n414 VGND.n413 54.0035
R768 VGND.n416 VGND.n412 54.0035
R769 VGND.n461 VGND.n379 53.9218
R770 VGND.n401 VGND.n400 53.9218
R771 VGND.n616 VGND.n615 53.3664
R772 VGND.n619 VGND.n618 53.3664
R773 VGND.n622 VGND.n621 53.3664
R774 VGND.n671 VGND.n545 53.3664
R775 VGND.n665 VGND.n547 53.3664
R776 VGND.n658 VGND.n549 53.3664
R777 VGND.n651 VGND.n552 53.3664
R778 VGND.n644 VGND.n555 53.3664
R779 VGND.n568 VGND.n567 53.3664
R780 VGND.n684 VGND.n683 53.3664
R781 VGND.n687 VGND.n686 53.3664
R782 VGND.n722 VGND.n263 53.3664
R783 VGND.n720 VGND.n719 53.3664
R784 VGND.n711 VGND.n271 53.3664
R785 VGND.n709 VGND.n708 53.3664
R786 VGND.n146 VGND.n28 53.3664
R787 VGND.n79 VGND.n29 53.3664
R788 VGND.n135 VGND.n30 53.3664
R789 VGND.n129 VGND.n31 53.3664
R790 VGND.n147 VGND.n26 53.3664
R791 VGND.n150 VGND.n33 53.3664
R792 VGND.n164 VGND.n35 53.3664
R793 VGND.n176 VGND.n40 53.3664
R794 VGND.n194 VGND.n44 53.3664
R795 VGND.n204 VGND.n43 53.3664
R796 VGND.n208 VGND.n42 53.3664
R797 VGND.n217 VGND.n41 53.3664
R798 VGND.n110 VGND.n27 53.3664
R799 VGND.n105 VGND.n34 53.3664
R800 VGND.n38 VGND.n37 53.3664
R801 VGND.n775 VGND.n774 53.3664
R802 VGND.n774 VGND.n25 53.3664
R803 VGND.n38 VGND.n24 53.3664
R804 VGND.n36 VGND.n34 53.3664
R805 VGND.n106 VGND.n27 53.3664
R806 VGND.n78 VGND.n28 53.3664
R807 VGND.n136 VGND.n29 53.3664
R808 VGND.n130 VGND.n30 53.3664
R809 VGND.n123 VGND.n31 53.3664
R810 VGND.n45 VGND.n40 53.3664
R811 VGND.n167 VGND.n35 53.3664
R812 VGND.n163 VGND.n33 53.3664
R813 VGND.n151 VGND.n26 53.3664
R814 VGND.n207 VGND.n41 53.3664
R815 VGND.n205 VGND.n42 53.3664
R816 VGND.n193 VGND.n43 53.3664
R817 VGND.n46 VGND.n44 53.3664
R818 VGND.n710 VGND.n709 53.3664
R819 VGND.n271 VGND.n265 53.3664
R820 VGND.n721 VGND.n720 53.3664
R821 VGND.n592 VGND.n263 53.3664
R822 VGND.n623 VGND.n622 53.3664
R823 VGND.n620 VGND.n619 53.3664
R824 VGND.n617 VGND.n616 53.3664
R825 VGND.n666 VGND.n545 53.3664
R826 VGND.n659 VGND.n547 53.3664
R827 VGND.n652 VGND.n549 53.3664
R828 VGND.n645 VGND.n552 53.3664
R829 VGND.n688 VGND.n687 53.3664
R830 VGND.n685 VGND.n684 53.3664
R831 VGND.n567 VGND.n292 53.3664
R832 VGND.n566 VGND.n555 53.3664
R833 VGND.n444 VGND.n394 53.1823
R834 VGND.n444 VGND.t56 53.1823
R835 VGND.n428 VGND.n392 53.1823
R836 VGND.t56 VGND.n392 53.1823
R837 VGND.n302 VGND.n300 53.1823
R838 VGND.n300 VGND.t54 53.1823
R839 VGND.n301 VGND.n299 53.1823
R840 VGND.n299 VGND.t54 53.1823
R841 VGND.n472 VGND.n471 48.7505
R842 VGND.n471 VGND.n470 48.7505
R843 VGND.n353 VGND.n352 48.7505
R844 VGND.n354 VGND.n353 48.7505
R845 VGND.n430 VGND.n429 42.0571
R846 VGND.n506 VGND.n505 42.0571
R847 VGND.n428 VGND.n390 41.1681
R848 VGND.n306 VGND.n301 41.1681
R849 VGND.n454 VGND.n384 39.7638
R850 VGND.n457 VGND.n456 39.511
R851 VGND.n469 VGND.n335 36.4578
R852 VGND.t11 VGND.t38 35.1962
R853 VGND.t18 VGND.t19 35.1962
R854 VGND.t39 VGND.t24 35.1962
R855 VGND.t26 VGND.t10 35.1962
R856 VGND.n429 VGND.n393 34.4123
R857 VGND.n443 VGND.n393 34.4123
R858 VGND.n446 VGND.n445 34.4123
R859 VGND.n445 VGND.n387 34.4123
R860 VGND.n507 VGND.n506 34.4123
R861 VGND.n508 VGND.n507 34.4123
R862 VGND.n501 VGND.n500 34.4123
R863 VGND.n500 VGND.n499 34.4123
R864 VGND.n489 VGND.n313 34.4123
R865 VGND.t40 VGND.n313 34.4123
R866 VGND.n368 VGND.n312 34.4123
R867 VGND.t40 VGND.n312 34.4123
R868 VGND.n466 VGND.n332 33.9329
R869 VGND.n450 VGND.t33 33.4483
R870 VGND.n334 VGND.n331 32.5005
R871 VGND.t58 VGND.n334 32.5005
R872 VGND.n333 VGND.n319 32.5005
R873 VGND.t58 VGND.n333 32.5005
R874 VGND.n454 VGND.n453 32.5005
R875 VGND.n453 VGND.n452 32.5005
R876 VGND.n410 VGND.n409 32.5005
R877 VGND.n409 VGND.n408 32.5005
R878 VGND.n530 VGND.n296 32.4888
R879 VGND.t40 VGND.n361 32.28
R880 VGND.n47 VGND.n4 32.1396
R881 VGND.n756 VGND.n755 32.1396
R882 VGND.n394 VGND.t57 30.8834
R883 VGND.n302 VGND.t55 30.8834
R884 VGND.n371 VGND.n370 30.4707
R885 VGND.n361 VGND.n360 28.2867
R886 VGND.n347 VGND.n331 28.0594
R887 VGND.n679 VGND.t82 26.9203
R888 VGND.n527 VGND.t24 26.8034
R889 VGND.n574 VGND.t86 26.6016
R890 VGND.n795 VGND.t7 26.5326
R891 VGND.n790 VGND.t22 26.5035
R892 VGND.t19 VGND.n509 25.9911
R893 VGND.n239 VGND.t4 25.1357
R894 VGND.n12 VGND.t51 25.0376
R895 VGND.n485 VGND.n484 24.7516
R896 VGND.t82 VGND.n588 24.6974
R897 VGND.n337 VGND.n332 24.4644
R898 VGND.n297 VGND.t7 23.9031
R899 VGND.n510 VGND.t11 23.8874
R900 VGND.n575 VGND.n244 23.8095
R901 VGND.n516 VGND.n8 23.4151
R902 VGND.n739 VGND.n737 23.4151
R903 VGND.n434 VGND.n433 23.0405
R904 VGND.n503 VGND.n303 23.0405
R905 VGND.t63 VGND.t40 22.9622
R906 VGND.n520 VGND.n519 22.5696
R907 VGND.n607 VGND.n247 21.7338
R908 VGND.n802 VGND.n801 21.6664
R909 VGND.n296 VGND.n232 20.8472
R910 VGND.n580 VGND.n571 20.7857
R911 VGND.n579 VGND.n572 20.7857
R912 VGND.n574 VGND.n573 20.7857
R913 VGND.n398 VGND.n397 20.7665
R914 VGND.n243 VGND.n242 20.7665
R915 VGND.n750 VGND.n241 20.7665
R916 VGND.n751 VGND.n240 20.7665
R917 VGND.n790 VGND.n789 20.6876
R918 VGND.n788 VGND.n10 20.6876
R919 VGND.n787 VGND.n11 20.6876
R920 VGND.n2 VGND.n1 20.6683
R921 VGND.n799 VGND.n798 20.6683
R922 VGND.n802 VGND.n800 20.6683
R923 VGND.n490 VGND.n314 20.517
R924 VGND.n492 VGND.n311 20.3
R925 VGND.n338 VGND.n337 20.1729
R926 VGND.n345 VGND.n338 20.1729
R927 VGND.n375 VGND.n336 20.1729
R928 VGND.n345 VGND.n336 20.1729
R929 VGND.n362 VGND.n314 20.0772
R930 VGND.n475 VGND.n474 19.4026
R931 VGND.n351 VGND.n347 19.2005
R932 VGND.n468 VGND.n467 18.8715
R933 VGND.n469 VGND.n468 18.8715
R934 VGND.n356 VGND.n355 18.8715
R935 VGND.n357 VGND.n356 18.8715
R936 VGND.n451 VGND.n231 18.7538
R937 VGND.n446 VGND.n391 18.7337
R938 VGND.n502 VGND.n501 18.7337
R939 VGND.n737 VGND.n252 17.5097
R940 VGND.n792 VGND.n9 17.2467
R941 VGND.n485 VGND.n318 17.1218
R942 VGND.n474 VGND.n473 16.4046
R943 VGND.n447 VGND.n446 16.3845
R944 VGND.n501 VGND.n304 16.3845
R945 VGND.n793 VGND.n8 16.2573
R946 VGND.n472 VGND.n332 16.1396
R947 VGND.n577 VGND.n576 16.0068
R948 VGND.n420 VGND.n419 15.5385
R949 VGND.n47 VGND.n6 14.6255
R950 VGND.n762 VGND.n6 14.6255
R951 VGND.n7 VGND.n5 14.6255
R952 VGND.n513 VGND.n7 14.6255
R953 VGND.n757 VGND.n756 14.6255
R954 VGND.n758 VGND.n757 14.6255
R955 VGND.n746 VGND.n745 14.6255
R956 VGND.n354 VGND.t77 14.0932
R957 VGND.n480 VGND.n323 14.0913
R958 VGND.n474 VGND.n326 12.7191
R959 VGND.n530 VGND.t10 12.4544
R960 VGND.n448 VGND.n447 11.9393
R961 VGND.n449 VGND.n448 11.9393
R962 VGND.n436 VGND.n435 11.9393
R963 VGND.n437 VGND.n436 11.9393
R964 VGND.n497 VGND.n304 11.9393
R965 VGND.n498 VGND.n497 11.9393
R966 VGND.n309 VGND.n308 11.9393
R967 VGND.n494 VGND.n309 11.9393
R968 VGND.t16 VGND.n743 11.7213
R969 VGND.n379 VGND.t76 11.6005
R970 VGND.n379 VGND.t79 11.6005
R971 VGND.n400 VGND.t74 11.6005
R972 VGND.n400 VGND.t75 11.6005
R973 VGND.n413 VGND.t80 11.6005
R974 VGND.n413 VGND.t68 11.6005
R975 VGND.n412 VGND.t70 11.6005
R976 VGND.n412 VGND.t72 11.6005
R977 VGND.n458 VGND.n381 10.5495
R978 VGND.t39 VGND.n510 10.2545
R979 VGND.n394 VGND.n391 10.0532
R980 VGND.n502 VGND.n302 10.0532
R981 VGND.n371 VGND.n316 9.74099
R982 VGND.n439 VGND.n438 9.6713
R983 VGND.n141 VGND.n71 9.36638
R984 VGND.n346 VGND.n327 9.3005
R985 VGND.n457 VGND.n380 9.3005
R986 VGND.n422 VGND.n421 9.3005
R987 VGND.n423 VGND.n383 9.3005
R988 VGND.n367 VGND.n314 8.86924
R989 VGND.t38 VGND.n509 8.66405
R990 VGND.n795 VGND.t27 8.66405
R991 VGND.n488 VGND.n315 8.42977
R992 VGND.n527 VGND.t27 7.85184
R993 VGND.n434 VGND.n389 7.5005
R994 VGND.n395 VGND.n389 7.5005
R995 VGND.n396 VGND.n388 7.5005
R996 VGND.n395 VGND.n388 7.5005
R997 VGND.n496 VGND.n303 7.5005
R998 VGND.n496 VGND.n495 7.5005
R999 VGND.n307 VGND.n305 7.5005
R1000 VGND.n495 VGND.n305 7.5005
R1001 VGND.n484 VGND.n319 7.34725
R1002 VGND.n487 VGND.n486 7.32557
R1003 VGND.n519 VGND.n518 7.313
R1004 VGND.n518 VGND.n517 7.313
R1005 VGND.n523 VGND.n522 7.313
R1006 VGND.n524 VGND.n523 7.313
R1007 VGND.n575 VGND.n251 7.313
R1008 VGND.n588 VGND.n251 7.313
R1009 VGND.n740 VGND.n250 7.313
R1010 VGND.n604 VGND.n250 7.313
R1011 VGND.t18 VGND.n514 7.03963
R1012 VGND.n486 VGND.n485 6.9983
R1013 VGND.n806 VGND.n805 6.9005
R1014 VGND.n4 VGND.n3 6.9005
R1015 VGND.n755 VGND.n754 6.9005
R1016 VGND.n753 VGND.n238 6.9005
R1017 VGND.n328 VGND 6.21282
R1018 VGND.n797 VGND.n796 6.15839
R1019 VGND.n796 VGND.n795 6.15839
R1020 VGND.n794 VGND.n793 6.15839
R1021 VGND.n795 VGND.n794 6.15839
R1022 VGND.n747 VGND.n236 6.15839
R1023 VGND.n236 VGND.n235 6.15839
R1024 VGND.n252 VGND.n234 6.15839
R1025 VGND.n246 VGND.n234 6.15839
R1026 VGND.n370 VGND.n369 5.92892
R1027 VGND.n487 VGND.n316 5.77749
R1028 VGND.n368 VGND.n367 5.73359
R1029 VGND.t58 VGND.n345 5.51505
R1030 VGND.n370 VGND.n342 5.34506
R1031 VGND.n425 VGND 5.06219
R1032 VGND.t16 VGND.n247 4.93988
R1033 VGND.n118 VGND.n87 4.90263
R1034 VGND.n91 VGND.n66 4.90263
R1035 VGND.n599 VGND.n542 4.90263
R1036 VGND.n561 VGND.n556 4.90263
R1037 VGND.n386 VGND.n381 4.8755
R1038 VGND.n438 VGND.n386 4.8755
R1039 VGND.n419 VGND.n385 4.8755
R1040 VGND.n438 VGND.n385 4.8755
R1041 VGND.n148 VGND.n66 4.84816
R1042 VGND.n153 VGND.n152 4.84816
R1043 VGND.n149 VGND.n62 4.84816
R1044 VGND.n165 VGND.n61 4.84816
R1045 VGND.n169 VGND.n168 4.84816
R1046 VGND.n166 VGND.n58 4.84816
R1047 VGND.n177 VGND.n175 4.84816
R1048 VGND.n179 VGND.n178 4.84816
R1049 VGND.n643 VGND.n556 4.84816
R1050 VGND.n642 VGND.n557 4.84816
R1051 VGND.n569 VGND.n565 4.84816
R1052 VGND.n682 VGND.n293 4.84816
R1053 VGND.n681 VGND.n291 4.84816
R1054 VGND.n290 VGND.n286 4.84816
R1055 VGND.n690 VGND.n689 4.84816
R1056 VGND.n287 VGND.n282 4.84816
R1057 VGND.n765 VGND.n54 4.57193
R1058 VGND.n700 VGND.n281 4.57193
R1059 VGND.n403 VGND.n380 4.5005
R1060 VGND.n328 VGND.n326 4.5005
R1061 VGND.n464 VGND.n322 4.5005
R1062 VGND.n348 VGND.n327 4.5005
R1063 VGND.n422 VGND.n406 4.5005
R1064 VGND.n424 VGND.n423 4.5005
R1065 VGND.n397 VGND.t15 4.3505
R1066 VGND.n397 VGND.t14 4.3505
R1067 VGND.n242 VGND.t20 4.3505
R1068 VGND.n242 VGND.t9 4.3505
R1069 VGND.n241 VGND.t23 4.3505
R1070 VGND.n241 VGND.t29 4.3505
R1071 VGND.n240 VGND.t31 4.3505
R1072 VGND.n240 VGND.t52 4.3505
R1073 VGND.n789 VGND.t2 4.3505
R1074 VGND.n789 VGND.t41 4.3505
R1075 VGND.n10 VGND.t32 4.3505
R1076 VGND.n10 VGND.t50 4.3505
R1077 VGND.n11 VGND.t85 4.3505
R1078 VGND.n11 VGND.t36 4.3505
R1079 VGND.n1 VGND.t37 4.3505
R1080 VGND.n1 VGND.t42 4.3505
R1081 VGND.n798 VGND.t47 4.3505
R1082 VGND.n798 VGND.t49 4.3505
R1083 VGND.n800 VGND.t44 4.3505
R1084 VGND.n800 VGND.t88 4.3505
R1085 VGND.n801 VGND.t53 4.3505
R1086 VGND.n801 VGND.t12 4.3505
R1087 VGND.n571 VGND.t87 4.3505
R1088 VGND.n571 VGND.t61 4.3505
R1089 VGND.n572 VGND.t46 4.3505
R1090 VGND.n572 VGND.t28 4.3505
R1091 VGND.n573 VGND.t25 4.3505
R1092 VGND.n573 VGND.t45 4.3505
R1093 VGND.n809 VGND 4.3492
R1094 VGND.n432 VGND.n424 4.26937
R1095 VGND.n417 VGND.n411 4.25229
R1096 VGND.n422 VGND.n407 4.1668
R1097 VGND.n12 VGND.n3 4.10351
R1098 VGND.n754 VGND.n239 4.10351
R1099 VGND.n232 VGND.t5 4.05043
R1100 VGND.n417 VGND.n416 4.02718
R1101 VGND.n355 VGND.n317 3.98739
R1102 VGND.n767 VGND.n48 3.9624
R1103 VGND.n279 VGND.n237 3.9624
R1104 VGND.n629 VGND.n588 3.952
R1105 VGND.t39 VGND.n511 3.92193
R1106 VGND.n98 VGND.n87 3.81327
R1107 VGND.n112 VGND.n111 3.81327
R1108 VGND.n108 VGND.n107 3.81327
R1109 VGND.n104 VGND.n102 3.81327
R1110 VGND.n103 VGND.n15 3.81327
R1111 VGND.n783 VGND.n16 3.81327
R1112 VGND.n22 VGND.n21 3.81327
R1113 VGND.n777 VGND.n776 3.81327
R1114 VGND.n220 VGND.n23 3.81327
R1115 VGND.n601 VGND.n599 3.81327
R1116 VGND.n603 VGND.n602 3.81327
R1117 VGND.n614 VGND.n597 3.81327
R1118 VGND.n613 VGND.n595 3.81327
R1119 VGND.n594 VGND.n584 3.81327
R1120 VGND.n631 VGND.n585 3.81327
R1121 VGND.n590 VGND.n589 3.81327
R1122 VGND.n625 VGND.n624 3.81327
R1123 VGND.n591 VGND.n255 3.81327
R1124 VGND.n421 VGND.n384 3.76521
R1125 VGND.n430 VGND.n394 3.71562
R1126 VGND.n505 VGND.n302 3.71562
R1127 VGND.n54 VGND.n53 3.55606
R1128 VGND.n698 VGND.n281 3.55606
R1129 VGND.n297 VGND.t26 3.54046
R1130 VGND.n162 VGND.n161 3.48646
R1131 VGND.n635 VGND.n570 3.48646
R1132 VGND.n504 VGND.n503 3.46869
R1133 VGND.n432 VGND.n431 3.33015
R1134 VGND.n323 VGND.t59 3.16414
R1135 VGND.n323 VGND.t60 3.16414
R1136 VGND.n418 VGND.n417 3.10035
R1137 VGND.n475 VGND.n331 2.96471
R1138 VGND.n426 VGND 2.88148
R1139 VGND.n145 VGND.n144 2.7239
R1140 VGND.n77 VGND.n68 2.7239
R1141 VGND.n138 VGND.n80 2.7239
R1142 VGND.n134 VGND.n133 2.7239
R1143 VGND.n131 VGND.n83 2.7239
R1144 VGND.n128 VGND.n127 2.7239
R1145 VGND.n124 VGND.n85 2.7239
R1146 VGND.n121 VGND.n120 2.7239
R1147 VGND.n674 VGND.n673 2.7239
R1148 VGND.n670 VGND.n543 2.7239
R1149 VGND.n669 VGND.n667 2.7239
R1150 VGND.n664 VGND.n546 2.7239
R1151 VGND.n663 VGND.n660 2.7239
R1152 VGND.n656 VGND.n653 2.7239
R1153 VGND.n650 VGND.n551 2.7239
R1154 VGND.n649 VGND.n646 2.7239
R1155 VGND.n376 VGND.n374 2.68591
R1156 VGND VGND.n0 2.56118
R1157 VGND.n462 VGND.n461 2.53642
R1158 VGND.n372 VGND.n371 2.3255
R1159 VGND.n459 VGND.n380 2.29617
R1160 VGND.n806 VGND.n3 2.28754
R1161 VGND.n754 VGND.n753 2.28754
R1162 VGND.n145 VGND.n67 2.17922
R1163 VGND.n144 VGND.n68 2.17922
R1164 VGND.n80 VGND.n77 2.17922
R1165 VGND.n138 VGND.n137 2.17922
R1166 VGND.n134 VGND.n82 2.17922
R1167 VGND.n133 VGND.n131 2.17922
R1168 VGND.n128 VGND.n83 2.17922
R1169 VGND.n127 VGND.n124 2.17922
R1170 VGND.n121 VGND.n85 2.17922
R1171 VGND.n673 VGND.n543 2.17922
R1172 VGND.n670 VGND.n669 2.17922
R1173 VGND.n667 VGND.n546 2.17922
R1174 VGND.n664 VGND.n663 2.17922
R1175 VGND.n660 VGND.n548 2.17922
R1176 VGND.n657 VGND.n656 2.17922
R1177 VGND.n653 VGND.n551 2.17922
R1178 VGND.n650 VGND.n649 2.17922
R1179 VGND.n646 VGND.n554 2.17922
R1180 VGND.n227 VGND.n219 2.17819
R1181 VGND.n259 VGND.n254 2.17819
R1182 VGND.n416 VGND.n415 2.15904
R1183 VGND.n414 VGND.n406 2.12067
R1184 VGND.n377 VGND.n376 2.10102
R1185 VGND.n426 VGND.n425 2.08765
R1186 VGND.n192 VGND.n13 1.89157
R1187 VGND.n582 VGND.n581 1.89157
R1188 VGND.n470 VGND.t78 1.83868
R1189 VGND.n771 VGND.n49 1.79105
R1190 VGND.n196 VGND.n190 1.79105
R1191 VGND.n203 VGND.n201 1.79105
R1192 VGND.n210 VGND.n209 1.79105
R1193 VGND.n188 VGND.n187 1.79105
R1194 VGND.n218 VGND.n216 1.79105
R1195 VGND.n724 VGND.n261 1.79105
R1196 VGND.n723 VGND.n262 1.79105
R1197 VGND.n266 VGND.n264 1.79105
R1198 VGND.n718 VGND.n717 1.79105
R1199 VGND.n713 VGND.n267 1.79105
R1200 VGND.n707 VGND.n706 1.79105
R1201 VGND.n415 VGND.n414 1.78099
R1202 VGND.n206 VGND 1.76685
R1203 VGND.n505 VGND.n504 1.7255
R1204 VGND.n431 VGND.n430 1.7255
R1205 VGND.n9 VGND 1.71609
R1206 VGND.n576 VGND 1.7155
R1207 VGND.n399 VGND.n0 1.71444
R1208 VGND.n550 VGND.n548 1.68901
R1209 VGND.n736 VGND.n735 1.64587
R1210 VGND.n82 VGND.n81 1.63454
R1211 VGND.n226 VGND.n225 1.62167
R1212 VGND.n810 VGND.n0 1.58664
R1213 VGND.n374 VGND.n373 1.55732
R1214 VGND.n161 VGND.n14 1.51978
R1215 VGND.n635 VGND.n634 1.51978
R1216 VGND.n525 VGND.n511 1.4937
R1217 VGND.n369 VGND.n368 1.47378
R1218 VGND.n788 VGND.n787 1.46641
R1219 VGND.n580 VGND.n579 1.46641
R1220 VGND.n578 VGND.n574 1.43989
R1221 VGND.n791 VGND.n790 1.43895
R1222 VGND.n463 VGND.n462 1.43287
R1223 VGND.n810 VGND.n809 1.42519
R1224 VGND VGND.n427 1.412
R1225 VGND.n772 VGND.n48 1.37971
R1226 VGND.n272 VGND 1.37971
R1227 VGND.n276 VGND.n237 1.37971
R1228 VGND.n161 VGND.n160 1.3622
R1229 VGND.n636 VGND.n635 1.3622
R1230 VGND.n456 VGND.n455 1.30961
R1231 VGND.n402 VGND.n399 1.30876
R1232 VGND.n425 VGND 1.24253
R1233 VGND.n192 VGND.n191 1.21033
R1234 VGND.n461 VGND.n460 1.20454
R1235 VGND.n581 VGND.n275 1.18613
R1236 VGND.n767 VGND.n766 1.11796
R1237 VGND.n699 VGND.n279 1.11796
R1238 VGND.n402 VGND.n401 1.1014
R1239 VGND.n112 VGND.n98 1.08986
R1240 VGND.n111 VGND.n108 1.08986
R1241 VGND.n107 VGND.n102 1.08986
R1242 VGND.n104 VGND.n103 1.08986
R1243 VGND.n21 VGND.n16 1.08986
R1244 VGND.n777 VGND.n22 1.08986
R1245 VGND.n776 VGND.n23 1.08986
R1246 VGND.n224 VGND.n220 1.08986
R1247 VGND.n226 VGND.n224 1.08986
R1248 VGND.n137 VGND.n81 1.08986
R1249 VGND.n180 VGND.n53 1.08986
R1250 VGND.n603 VGND.n601 1.08986
R1251 VGND.n602 VGND.n597 1.08986
R1252 VGND.n614 VGND.n613 1.08986
R1253 VGND.n595 VGND.n594 1.08986
R1254 VGND.n589 VGND.n585 1.08986
R1255 VGND.n625 VGND.n590 1.08986
R1256 VGND.n624 VGND.n591 1.08986
R1257 VGND.n734 VGND.n255 1.08986
R1258 VGND.n735 VGND.n734 1.08986
R1259 VGND.n698 VGND.n697 1.08986
R1260 VGND.n808 VGND 1.08385
R1261 VGND.t30 VGND.t35 1.07946
R1262 VGND.t62 VGND.t33 1.07946
R1263 VGND.n463 VGND.n322 1.07186
R1264 VGND.n455 VGND.n454 1.06085
R1265 VGND.n465 VGND.n464 1.05279
R1266 VGND.n657 VGND.n550 1.03539
R1267 VGND.n466 VGND.n465 1.03383
R1268 VGND.n462 VGND.n378 1.0271
R1269 VGND.n398 VGND.n243 0.998567
R1270 VGND.n799 VGND.n2 0.997923
R1271 VGND.n751 VGND.n750 0.997923
R1272 VGND.n604 VGND.n533 0.988376
R1273 VGND.n784 VGND.n15 0.871989
R1274 VGND.n632 VGND.n584 0.871989
R1275 VGND.n401 VGND.n378 0.837944
R1276 VGND.n227 VGND.n226 0.823184
R1277 VGND.n119 VGND.n118 0.817521
R1278 VGND.n91 VGND.n90 0.817521
R1279 VGND.n675 VGND.n542 0.817521
R1280 VGND.n561 VGND.n560 0.817521
R1281 VGND.n735 VGND.n254 0.798988
R1282 VGND.n347 VGND.n346 0.775237
R1283 VGND.n634 VGND.n633 0.765632
R1284 VGND.n785 VGND.n14 0.764974
R1285 VGND.n793 VGND.n792 0.751968
R1286 VGND.n577 VGND.n252 0.739443
R1287 VGND.n384 VGND.n383 0.684992
R1288 VGND.n337 VGND.n319 0.682157
R1289 VGND.n786 VGND.n785 0.653909
R1290 VGND.n633 VGND.n583 0.653909
R1291 VGND.n808 VGND.n807 0.636285
R1292 VGND.n752 VGND.n751 0.633876
R1293 VGND.n581 VGND.n273 0.605415
R1294 VGND.n81 VGND.n14 0.596304
R1295 VGND.n634 VGND.n550 0.596304
R1296 VGND.n785 VGND.n784 0.59175
R1297 VGND.n633 VGND.n632 0.59175
R1298 VGND.n195 VGND.n192 0.581218
R1299 VGND.n787 VGND.n786 0.539326
R1300 VGND.n583 VGND.n580 0.539326
R1301 VGND.n804 VGND.n797 0.532356
R1302 VGND.n748 VGND.n747 0.532356
R1303 VGND.n803 VGND.n802 0.528206
R1304 VGND.n749 VGND.n243 0.528206
R1305 VGND.n405 VGND.n404 0.494548
R1306 VGND.n476 VGND.n327 0.47062
R1307 VGND.n803 VGND.n799 0.469572
R1308 VGND.n750 VGND.n749 0.469572
R1309 VGND.n382 VGND.n380 0.469344
R1310 VGND.t13 VGND.t48 0.461668
R1311 VGND.t34 VGND.t43 0.461668
R1312 VGND.n348 VGND.n330 0.456098
R1313 VGND.n583 VGND.n582 0.452967
R1314 VGND.n786 VGND.n13 0.452516
R1315 VGND.n483 VGND.n482 0.452003
R1316 VGND.n465 VGND.n463 0.4505
R1317 VGND.n423 VGND.n382 0.441368
R1318 VGND.n712 VGND 0.411842
R1319 VGND VGND.n811 0.406951
R1320 VGND.n807 VGND.n2 0.403851
R1321 VGND.n349 VGND.n348 0.399345
R1322 VGND.n376 VGND.n375 0.391918
R1323 VGND.n772 VGND.n771 0.387646
R1324 VGND.n191 VGND.n49 0.387646
R1325 VGND.n196 VGND.n195 0.387646
R1326 VGND.n201 VGND.n190 0.387646
R1327 VGND.n210 VGND.n206 0.387646
R1328 VGND.n209 VGND.n188 0.387646
R1329 VGND.n216 VGND.n187 0.387646
R1330 VGND.n219 VGND.n218 0.387646
R1331 VGND.n261 VGND.n259 0.387646
R1332 VGND.n724 VGND.n723 0.387646
R1333 VGND.n264 VGND.n262 0.387646
R1334 VGND.n718 VGND.n266 0.387646
R1335 VGND.n717 VGND.n267 0.387646
R1336 VGND.n273 VGND.n272 0.387646
R1337 VGND.n707 VGND.n275 0.387646
R1338 VGND.n706 VGND.n276 0.387646
R1339 VGND.n483 VGND.n320 0.376108
R1340 VGND.n807 VGND.n806 0.373405
R1341 VGND.n373 VGND.n372 0.368932
R1342 VGND.n372 VGND.n341 0.355
R1343 VGND.n477 VGND.n476 0.350102
R1344 VGND.n330 VGND.n329 0.344129
R1345 VGND.n753 VGND.n752 0.343093
R1346 VGND.n456 VGND.n382 0.32741
R1347 VGND.n120 VGND.n119 0.327309
R1348 VGND.n675 VGND.n674 0.327309
R1349 VGND.n482 VGND.n481 0.326722
R1350 VGND.n424 VGND.n405 0.317677
R1351 VGND.n349 VGND.n320 0.312188
R1352 VGND.n374 VGND.n317 0.3005
R1353 VGND.n350 VGND.n327 0.272145
R1354 VGND.n203 VGND 0.266663
R1355 VGND.n713 VGND 0.242466
R1356 VGND.n479 VGND.n324 0.226831
R1357 VGND.n352 VGND.n318 0.224276
R1358 VGND.n351 VGND.n350 0.221929
R1359 VGND.n482 VGND.n321 0.221128
R1360 VGND.n478 VGND.n477 0.220839
R1361 VGND.n784 VGND.n783 0.218372
R1362 VGND.n632 VGND.n631 0.218372
R1363 VGND.n481 VGND.n480 0.216846
R1364 VGND.n325 VGND.n321 0.20954
R1365 VGND.n811 VGND.n810 0.19179
R1366 VGND.n576 VGND.n575 0.188367
R1367 VGND.n316 VGND.n315 0.187817
R1368 VGND.n375 VGND.n339 0.180782
R1369 VGND.n519 VGND.n9 0.175842
R1370 VGND VGND.n712 0.14568
R1371 VGND.n433 VGND.n432 0.139042
R1372 VGND.n809 VGND.n808 0.135155
R1373 VGND.n473 VGND.n325 0.133357
R1374 VGND.n460 VGND.n378 0.131666
R1375 VGND.n484 VGND.n483 0.126176
R1376 VGND.n405 VGND.n382 0.1255
R1377 VGND.n369 VGND.n341 0.122868
R1378 VGND.n399 VGND.n398 0.122278
R1379 VGND VGND.n202 0.121483
R1380 VGND.n504 VGND 0.120187
R1381 VGND.n431 VGND 0.120187
R1382 VGND.n341 VGND.n340 0.118284
R1383 VGND.n90 VGND.n67 0.109436
R1384 VGND.n560 VGND.n554 0.109436
R1385 VGND.n476 VGND.n475 0.107397
R1386 VGND.n792 VGND.n791 0.0987955
R1387 VGND.n578 VGND.n577 0.0987955
R1388 VGND.n13 VGND.n12 0.0952653
R1389 VGND.n582 VGND.n239 0.0948141
R1390 VGND.n420 VGND.n407 0.0850455
R1391 VGND.n752 VGND 0.0849072
R1392 VGND.n403 VGND.n402 0.0828991
R1393 VGND.n404 VGND 0.0780908
R1394 VGND.n804 VGND.n803 0.0736577
R1395 VGND.n749 VGND.n748 0.0736577
R1396 VGND.n423 VGND.n422 0.0711522
R1397 VGND.n479 VGND.n478 0.0605
R1398 VGND.n807 VGND 0.057201
R1399 VGND.n153 VGND.n148 0.0549681
R1400 VGND.n152 VGND.n149 0.0549681
R1401 VGND.n160 VGND.n62 0.0549681
R1402 VGND.n162 VGND.n61 0.0549681
R1403 VGND.n169 VGND.n165 0.0549681
R1404 VGND.n168 VGND.n166 0.0549681
R1405 VGND.n175 VGND.n58 0.0549681
R1406 VGND.n178 VGND.n177 0.0549681
R1407 VGND.n180 VGND.n179 0.0549681
R1408 VGND.n643 VGND.n642 0.0549681
R1409 VGND.n565 VGND.n557 0.0549681
R1410 VGND.n636 VGND.n569 0.0549681
R1411 VGND.n570 VGND.n293 0.0549681
R1412 VGND.n682 VGND.n681 0.0549681
R1413 VGND.n291 VGND.n290 0.0549681
R1414 VGND.n690 VGND.n286 0.0549681
R1415 VGND.n689 VGND.n287 0.0549681
R1416 VGND.n697 VGND.n282 0.0549681
R1417 VGND.n766 VGND.n765 0.0512937
R1418 VGND.n700 VGND.n699 0.0512937
R1419 VGND VGND.n324 0.048119
R1420 VGND.n476 VGND.n330 0.0459545
R1421 VGND.n352 VGND.n351 0.0452552
R1422 VGND.n329 VGND.n328 0.0448787
R1423 VGND.n477 VGND.n326 0.0428729
R1424 VGND.n373 VGND.n320 0.0382747
R1425 VGND.n415 VGND.n411 0.0367903
R1426 VGND.n481 VGND.n322 0.0330444
R1427 VGND.n464 VGND.n321 0.0294548
R1428 VGND.n459 VGND.n458 0.0286818
R1429 VGND.n791 VGND.n788 0.0279621
R1430 VGND.n579 VGND.n578 0.0270152
R1431 VGND.n473 VGND.n472 0.027001
R1432 VGND.n404 VGND.n403 0.0268453
R1433 VGND.n525 VGND.n510 0.0250793
R1434 VGND.n202 VGND 0.0246966
R1435 VGND.n424 VGND.n406 0.0246098
R1436 VGND.n411 VGND.n407 0.0135435
R1437 VGND.n460 VGND.n459 0.0126951
R1438 VGND.n350 VGND.n349 0.00969913
R1439 VGND.n329 VGND.n324 0.00493787
R1440 VGND.n427 VGND.n426 0.00387038
R1441 VGND.n811 VGND 0.00366816
R1442 VGND.n480 VGND.n479 0.00234911
R1443 VGND.n478 VGND.n325 0.00191243
R1444 VGND.n533 VGND.n532 0.00101101
R1445 VGND.n427 VGND 0.000702223
R1446 ua[2].n0 ua[2].t2 21.6012
R1447 ua[2].n1 ua[2].t3 21.6012
R1448 ua[2] ua[2].n2 9.84984
R1449 ua[2].n1 ua[2].t0 8.85318
R1450 ua[2].n0 ua[2].t1 8.85318
R1451 ua[2] ua[2].n1 2.55816
R1452 ua[2] ua[2].n0 2.55816
R1453 ua[2].n2 ua[2] 1.2695
R1454 ua[2].n2 ua[2] 1.10863
R1455 a_18163_10306.t0 a_18163_10306.t1 134.761
R1456 a_18163_10306.t0 a_18163_10306.t2 134.73
R1457 a_18163_10306.t4 a_18163_10306.n0 21.102
R1458 a_18163_10306.n0 a_18163_10306.t0 1.0135
R1459 a_18163_10306.t3 a_18163_10306.n0 18.8969
R1460 a_12378_15906.n40 a_12378_15906.t28 190.305
R1461 a_12378_15906.t28 a_12378_15906.n39 190.305
R1462 a_12378_15906.t26 a_12378_15906.n32 190.305
R1463 a_12378_15906.n38 a_12378_15906.t26 190.305
R1464 a_12378_15906.t10 a_12378_15906.n26 190.305
R1465 a_12378_15906.n27 a_12378_15906.t10 190.305
R1466 a_12378_15906.t24 a_12378_15906.n24 190.305
R1467 a_12378_15906.n28 a_12378_15906.t24 190.305
R1468 a_12378_15906.t22 a_12378_15906.n17 190.305
R1469 a_12378_15906.n18 a_12378_15906.t22 190.305
R1470 a_12378_15906.t16 a_12378_15906.n15 190.305
R1471 a_12378_15906.n81 a_12378_15906.t16 190.305
R1472 a_12378_15906.n78 a_12378_15906.t18 190.305
R1473 a_12378_15906.n22 a_12378_15906.t18 190.305
R1474 a_12378_15906.t12 a_12378_15906.n21 190.305
R1475 a_12378_15906.n75 a_12378_15906.t12 190.305
R1476 a_12378_15906.t36 a_12378_15906.n50 190.305
R1477 a_12378_15906.n14 a_12378_15906.t36 190.305
R1478 a_12378_15906.t32 a_12378_15906.n48 190.305
R1479 a_12378_15906.n51 a_12378_15906.t32 190.305
R1480 a_12378_15906.t30 a_12378_15906.n67 190.305
R1481 a_12378_15906.n71 a_12378_15906.t30 190.305
R1482 a_12378_15906.t14 a_12378_15906.n69 190.305
R1483 a_12378_15906.n70 a_12378_15906.t14 190.305
R1484 a_12378_15906.n62 a_12378_15906.t20 190.305
R1485 a_12378_15906.t20 a_12378_15906.n42 190.305
R1486 a_12378_15906.t8 a_12378_15906.n63 190.305
R1487 a_12378_15906.n64 a_12378_15906.t8 190.305
R1488 a_12378_15906.n19 a_12378_15906.t38 95.1811
R1489 a_12378_15906.n57 a_12378_15906.t34 95.1783
R1490 a_12378_15906.n36 a_12378_15906.n35 22.3176
R1491 a_12378_15906.n46 a_12378_15906.n45 22.2301
R1492 a_12378_15906.n0 a_12378_15906.n83 22.2284
R1493 a_12378_15906.n8 a_12378_15906.n44 22.2284
R1494 a_12378_15906.n12 a_12378_15906.n53 22.2284
R1495 a_12378_15906.n55 a_12378_15906.n54 22.2284
R1496 a_12378_15906.n10 a_12378_15906.n60 22.2284
R1497 a_12378_15906.n59 a_12378_15906.n58 22.2284
R1498 a_12378_15906.n84 a_12378_15906.n4 22.2284
R1499 a_12378_15906.n5 a_12378_15906.n23 22.1884
R1500 a_12378_15906.n9 a_12378_15906.n30 22.1884
R1501 a_12378_15906.n1 a_12378_15906.n31 22.1884
R1502 a_12378_15906.n3 a_12378_15906.n74 22.1884
R1503 a_12378_15906.n2 a_12378_15906.n73 22.1884
R1504 a_12378_15906.n11 a_12378_15906.n33 22.1884
R1505 a_12378_15906.n7 a_12378_15906.n34 22.1884
R1506 a_12378_15906.n57 a_12378_15906.n41 11.5566
R1507 a_12378_15906.n20 a_12378_15906.n19 10.9335
R1508 a_12378_15906.n79 a_12378_15906.n78 9.89233
R1509 a_12378_15906.n67 a_12378_15906.n66 9.89233
R1510 a_12378_15906.n26 a_12378_15906.n20 9.80925
R1511 a_12378_15906.n41 a_12378_15906.n40 9.80925
R1512 a_12378_15906.n65 a_12378_15906.n64 9.48127
R1513 a_12378_15906.n14 a_12378_15906.n13 9.40378
R1514 a_12378_15906.n81 a_12378_15906.n80 9.39819
R1515 a_12378_15906.n59 a_12378_15906.n57 4.9275
R1516 a_12378_15906.n19 a_12378_15906.n4 4.79654
R1517 a_12378_15906.n7 a_12378_15906.n6 4.5005
R1518 a_12378_15906.n37 a_12378_15906.n36 4.5005
R1519 a_12378_15906.n68 a_12378_15906.n11 4.5005
R1520 a_12378_15906.n2 a_12378_15906.n72 4.5005
R1521 a_12378_15906.n3 a_12378_15906.n76 4.5005
R1522 a_12378_15906.n77 a_12378_15906.n1 4.5005
R1523 a_12378_15906.n25 a_12378_15906.n5 4.5005
R1524 a_12378_15906.n9 a_12378_15906.n29 4.5005
R1525 a_12378_15906.n61 a_12378_15906.n10 4.5005
R1526 a_12378_15906.n56 a_12378_15906.n43 4.5005
R1527 a_12378_15906.n12 a_12378_15906.n52 4.5005
R1528 a_12378_15906.n49 a_12378_15906.n47 4.5005
R1529 a_12378_15906.n16 a_12378_15906.n8 4.5005
R1530 a_12378_15906.n0 a_12378_15906.n82 4.5005
R1531 a_12378_15906.n83 a_12378_15906.t7 4.3505
R1532 a_12378_15906.n83 a_12378_15906.t17 4.3505
R1533 a_12378_15906.n44 a_12378_15906.t23 4.3505
R1534 a_12378_15906.n44 a_12378_15906.t3 4.3505
R1535 a_12378_15906.n45 a_12378_15906.t1 4.3505
R1536 a_12378_15906.n45 a_12378_15906.t37 4.3505
R1537 a_12378_15906.n53 a_12378_15906.t33 4.3505
R1538 a_12378_15906.n53 a_12378_15906.t42 4.3505
R1539 a_12378_15906.n54 a_12378_15906.t44 4.3505
R1540 a_12378_15906.n54 a_12378_15906.t9 4.3505
R1541 a_12378_15906.n60 a_12378_15906.t21 4.3505
R1542 a_12378_15906.n60 a_12378_15906.t45 4.3505
R1543 a_12378_15906.n58 a_12378_15906.t5 4.3505
R1544 a_12378_15906.n58 a_12378_15906.t35 4.3505
R1545 a_12378_15906.n23 a_12378_15906.t6 4.3505
R1546 a_12378_15906.n23 a_12378_15906.t11 4.3505
R1547 a_12378_15906.n30 a_12378_15906.t25 4.3505
R1548 a_12378_15906.n30 a_12378_15906.t40 4.3505
R1549 a_12378_15906.n31 a_12378_15906.t2 4.3505
R1550 a_12378_15906.n31 a_12378_15906.t19 4.3505
R1551 a_12378_15906.n74 a_12378_15906.t13 4.3505
R1552 a_12378_15906.n74 a_12378_15906.t43 4.3505
R1553 a_12378_15906.n73 a_12378_15906.t0 4.3505
R1554 a_12378_15906.n73 a_12378_15906.t31 4.3505
R1555 a_12378_15906.n33 a_12378_15906.t15 4.3505
R1556 a_12378_15906.n33 a_12378_15906.t47 4.3505
R1557 a_12378_15906.n34 a_12378_15906.t4 4.3505
R1558 a_12378_15906.n34 a_12378_15906.t29 4.3505
R1559 a_12378_15906.n35 a_12378_15906.t27 4.3505
R1560 a_12378_15906.n35 a_12378_15906.t46 4.3505
R1561 a_12378_15906.t39 a_12378_15906.n84 4.3505
R1562 a_12378_15906.n84 a_12378_15906.t41 4.3505
R1563 a_12378_15906.n5 a_12378_15906.n4 2.55258
R1564 a_12378_15906.n80 a_12378_15906.n20 1.86108
R1565 a_12378_15906.n80 a_12378_15906.n79 1.86108
R1566 a_12378_15906.n79 a_12378_15906.n13 1.86108
R1567 a_12378_15906.n66 a_12378_15906.n13 1.86108
R1568 a_12378_15906.n66 a_12378_15906.n65 1.86108
R1569 a_12378_15906.n65 a_12378_15906.n41 1.86108
R1570 a_12378_15906.n4 a_12378_15906.n0 1.20675
R1571 a_12378_15906.n7 a_12378_15906.n11 1.0755
R1572 a_12378_15906.n3 a_12378_15906.n2 1.0755
R1573 a_12378_15906.n1 a_12378_15906.n9 1.0755
R1574 a_12378_15906.n46 a_12378_15906.n8 1.0755
R1575 a_12378_15906.n55 a_12378_15906.n12 1.0755
R1576 a_12378_15906.n10 a_12378_15906.n59 1.0755
R1577 a_12378_15906.n52 a_12378_15906.n48 0.759759
R1578 a_12378_15906.n50 a_12378_15906.n49 0.756673
R1579 a_12378_15906.n63 a_12378_15906.n43 0.702205
R1580 a_12378_15906.n62 a_12378_15906.n61 0.700784
R1581 a_12378_15906.n76 a_12378_15906.n75 0.669534
R1582 a_12378_15906.n72 a_12378_15906.n71 0.668114
R1583 a_12378_15906.n39 a_12378_15906.n6 0.666693
R1584 a_12378_15906.n77 a_12378_15906.n22 0.665273
R1585 a_12378_15906.n29 a_12378_15906.n28 0.662432
R1586 a_12378_15906.n27 a_12378_15906.n25 0.661011
R1587 a_12378_15906.n38 a_12378_15906.n37 0.659208
R1588 a_12378_15906.n49 a_12378_15906.n14 0.647608
R1589 a_12378_15906.n52 a_12378_15906.n51 0.645562
R1590 a_12378_15906.n26 a_12378_15906.n25 0.632599
R1591 a_12378_15906.n29 a_12378_15906.n24 0.631182
R1592 a_12378_15906.n70 a_12378_15906.n68 0.629532
R1593 a_12378_15906.n78 a_12378_15906.n77 0.628338
R1594 a_12378_15906.n40 a_12378_15906.n6 0.626917
R1595 a_12378_15906.n72 a_12378_15906.n67 0.625497
R1596 a_12378_15906.n76 a_12378_15906.n21 0.62408
R1597 a_12378_15906.n37 a_12378_15906.n32 0.619882
R1598 a_12378_15906.n69 a_12378_15906.n68 0.594586
R1599 a_12378_15906.n61 a_12378_15906.n42 0.59283
R1600 a_12378_15906.n64 a_12378_15906.n43 0.591408
R1601 a_12378_15906.n82 a_12378_15906.n15 0.580689
R1602 a_12378_15906.n17 a_12378_15906.n16 0.57833
R1603 a_12378_15906.n9 a_12378_15906.n5 0.538
R1604 a_12378_15906.n0 a_12378_15906.n8 0.538
R1605 a_12378_15906.n2 a_12378_15906.n11 0.537105
R1606 a_12378_15906.n1 a_12378_15906.n3 0.536664
R1607 a_12378_15906.n18 a_12378_15906.n16 0.495783
R1608 a_12378_15906.n82 a_12378_15906.n81 0.493424
R1609 a_12378_15906.n51 a_12378_15906.n14 0.488952
R1610 a_12378_15906.n50 a_12378_15906.n48 0.486913
R1611 a_12378_15906.n40 a_12378_15906.n32 0.476043
R1612 a_12378_15906.n39 a_12378_15906.n38 0.476043
R1613 a_12378_15906.n26 a_12378_15906.n24 0.459739
R1614 a_12378_15906.n28 a_12378_15906.n27 0.459739
R1615 a_12378_15906.n78 a_12378_15906.n21 0.459739
R1616 a_12378_15906.n75 a_12378_15906.n22 0.459739
R1617 a_12378_15906.n69 a_12378_15906.n67 0.459739
R1618 a_12378_15906.n71 a_12378_15906.n70 0.459739
R1619 a_12378_15906.n64 a_12378_15906.n42 0.451587
R1620 a_12378_15906.n63 a_12378_15906.n62 0.451587
R1621 a_12378_15906.n36 a_12378_15906.n7 0.408833
R1622 a_12378_15906.n81 a_12378_15906.n18 0.405391
R1623 a_12378_15906.n17 a_12378_15906.n15 0.405391
R1624 a_12378_15906.n12 a_12378_15906.n47 0.395292
R1625 a_12378_15906.n10 a_12378_15906.n56 0.395292
R1626 a_12378_15906.n47 a_12378_15906.n46 0.143208
R1627 a_12378_15906.n56 a_12378_15906.n55 0.143208
R1628 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 936.04
R1629 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 235.982
R1630 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 235.978
R1631 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 190.305
R1632 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 190.305
R1633 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 190.305
R1634 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 190.305
R1635 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 190.305
R1636 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 190.305
R1637 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 95.3928
R1638 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 95.3648
R1639 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 95.1789
R1640 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 95.1648
R1641 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 95.1542
R1642 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 95.1535
R1643 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 94.8314
R1644 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 94.8314
R1645 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 94.8314
R1646 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 94.8314
R1647 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 94.8314
R1648 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 94.8314
R1649 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 94.8314
R1650 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 94.8314
R1651 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 94.8314
R1652 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 94.8314
R1653 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 94.8314
R1654 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 94.8314
R1655 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 94.8314
R1656 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 94.8314
R1657 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 94.8314
R1658 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 94.8314
R1659 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 94.8314
R1660 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 94.8314
R1661 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 94.8314
R1662 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 94.8314
R1663 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 94.8314
R1664 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 94.8314
R1665 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 94.8314
R1666 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 84.0884
R1667 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 83.5719
R1668 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 83.5719
R1669 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 83.5719
R1670 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 83.5719
R1671 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 73.19
R1672 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 26.074
R1673 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 26.074
R1674 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 26.074
R1675 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 25.7843
R1676 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 10.2822
R1677 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 9.66398
R1678 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R1679 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R1680 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R1681 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R1682 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R1683 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 9.3005
R1684 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R1685 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R1686 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 9.3005
R1687 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R1688 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R1689 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R1690 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R1691 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R1692 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R1693 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R1694 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R1695 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R1696 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R1697 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R1698 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R1699 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R1700 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 9.3005
R1701 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R1702 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R1703 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 9.3005
R1704 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 9.3005
R1705 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 9.3005
R1706 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 7.22993
R1707 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 7.22993
R1708 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 7.22993
R1709 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 6.83022
R1710 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 6.81633
R1711 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 6.81633
R1712 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 6.81633
R1713 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 6.75312
R1714 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 4.64588
R1715 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 4.64588
R1716 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 4.64588
R1717 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 4.64588
R1718 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 2.29815
R1719 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 1.86108
R1720 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 1.86108
R1721 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 1.86108
R1722 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 1.86108
R1723 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 1.86108
R1724 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 1.86108
R1725 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 1.86108
R1726 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 1.28692
R1727 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 1.25468
R1728 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 1.14402
R1729 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 1.1424
R1730 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 1.12066
R1731 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 1.12066
R1732 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 1.11251
R1733 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 1.10979
R1734 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 1.10164
R1735 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 1.10164
R1736 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 1.10164
R1737 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 1.10164
R1738 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 1.09892
R1739 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 1.09349
R1740 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 1.09349
R1741 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 1.08805
R1742 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 1.08262
R1743 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 1.08262
R1744 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 1.08262
R1745 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 1.07024
R1746 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 1.0237
R1747 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.959578
R1748 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 0.812055
R1749 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.77514
R1750 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.701365
R1751 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.645119
R1752 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 0.645119
R1753 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 0.645119
R1754 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 0.645119
R1755 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 0.645119
R1756 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 0.645119
R1757 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 0.645119
R1758 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.645119
R1759 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 0.645119
R1760 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.645119
R1761 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 0.645119
R1762 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 0.645119
R1763 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 0.645119
R1764 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 0.645119
R1765 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 0.645119
R1766 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.645119
R1767 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 0.645119
R1768 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.645119
R1769 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 0.645119
R1770 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 0.645119
R1771 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 0.645119
R1772 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 0.645119
R1773 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 0.645119
R1774 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.645119
R1775 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.645119
R1776 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 0.645119
R1777 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 0.645119
R1778 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 0.645119
R1779 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 0.645119
R1780 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 0.645118
R1781 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 0.590702
R1782 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 0.572258
R1783 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 0.495065
R1784 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.495065
R1785 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 0.481478
R1786 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.481478
R1787 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.475521
R1788 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 0.470609
R1789 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.470609
R1790 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 0.465174
R1791 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 0.465174
R1792 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.465174
R1793 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.459844
R1794 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 0.459739
R1795 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.459739
R1796 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 0.446152
R1797 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.446152
R1798 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.445943
R1799 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.443435
R1800 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.440717
R1801 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 0.440717
R1802 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.434551
R1803 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 0.432263
R1804 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.414484
R1805 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.408265
R1806 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.408265
R1807 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.40372
R1808 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.40372
R1809 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.314045
R1810 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 0.290206
R1811 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.0183279
R1812 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 0.0112346
R1813 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 0.0112346
R1814 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 0.0112346
R1815 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 0.0112346
R1816 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.0112346
R1817 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 0.0112346
R1818 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 0.0112346
R1819 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 0.0112346
R1820 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 0.00759293
R1821 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 0.00316393
R1822 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t3 651.943
R1823 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t1 651.74
R1824 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t22 60.1752
R1825 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t25 60.1752
R1826 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t15 28.5589
R1827 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t10 27.6016
R1828 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n4 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t20 26.8562
R1829 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n4 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t26 26.0492
R1830 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n5 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t23 26.0492
R1831 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n6 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t24 26.0492
R1832 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n2 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t21 26.0492
R1833 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n10 24.2089
R1834 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n12 23.2516
R1835 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n11 23.2516
R1836 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n9 23.2516
R1837 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n8 23.2516
R1838 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n7 23.2516
R1839 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n13 23.2516
R1840 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t2 23
R1841 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t0 23
R1842 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n0 6.43084
R1843 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n12 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t8 4.3505
R1844 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n12 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t12 4.3505
R1845 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n11 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t19 4.3505
R1846 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n11 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t17 4.3505
R1847 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n10 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t11 4.3505
R1848 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n10 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t14 4.3505
R1849 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n9 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t9 4.3505
R1850 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n9 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t7 4.3505
R1851 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n8 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t5 4.3505
R1852 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n8 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t13 4.3505
R1853 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n7 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t18 4.3505
R1854 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n7 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t6 4.3505
R1855 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n13 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t16 4.3505
R1856 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n13 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t4 4.3505
R1857 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n1 3.89276
R1858 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n2 3.86689
R1859 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n5 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n4 2.80213
R1860 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n2 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n6 2.76952
R1861 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n6 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n5 2.72333
R1862 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t0 88.7532
R1863 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n14 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n12 22.2005
R1864 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n1 21.8665
R1865 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n16 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n15 21.5445
R1866 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n14 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n13 21.5445
R1867 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n20 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n19 21.5445
R1868 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n22 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n21 21.5445
R1869 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n24 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n23 21.5445
R1870 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n26 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n25 21.5445
R1871 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n29 21.5445
R1872 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n11 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n10 21.5445
R1873 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n9 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n8 21.5445
R1874 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n7 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n6 21.5445
R1875 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n5 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n4 21.5445
R1876 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n2 21.5445
R1877 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n18 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n17 21.5445
R1878 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n28 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n27 21.5418
R1879 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n15 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t19 4.3505
R1880 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n15 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t2 4.3505
R1881 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n13 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t4 4.3505
R1882 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n13 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t17 4.3505
R1883 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n12 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t26 4.3505
R1884 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n12 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t8 4.3505
R1885 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n19 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t20 4.3505
R1886 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n19 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t14 4.3505
R1887 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n21 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t15 4.3505
R1888 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n21 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t29 4.3505
R1889 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n23 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t18 4.3505
R1890 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n23 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t1 4.3505
R1891 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n25 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t5 4.3505
R1892 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n25 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t21 4.3505
R1893 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n27 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t30 4.3505
R1894 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n27 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t12 4.3505
R1895 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n29 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t9 4.3505
R1896 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n29 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t31 4.3505
R1897 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n10 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t25 4.3505
R1898 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n10 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t6 4.3505
R1899 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n8 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t3 4.3505
R1900 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n8 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t32 4.3505
R1901 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n6 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t23 4.3505
R1902 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n6 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t7 4.3505
R1903 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n4 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t10 4.3505
R1904 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n4 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t27 4.3505
R1905 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n2 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t28 4.3505
R1906 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n2 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t11 4.3505
R1907 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t13 4.3505
R1908 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t22 4.3505
R1909 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n17 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t16 4.3505
R1910 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n17 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t24 4.3505
R1911 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n28 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n26 1.51316
R1912 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n18 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n16 0.624699
R1913 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n26 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n24 0.624699
R1914 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n22 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n20 0.624699
R1915 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n5 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n3 0.60872
R1916 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n9 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n7 0.60872
R1917 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n11 0.553215
R1918 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n0 0.438342
R1919 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n0 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n28 0.298079
R1920 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n16 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n14 0.296969
R1921 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n24 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n22 0.296969
R1922 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n20 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n18 0.296969
R1923 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n7 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n5 0.289615
R1924 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n11 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n9 0.289615
R1925 VDPWR.n215 VDPWR.n104 17565.9
R1926 VDPWR.n217 VDPWR.n104 17565.9
R1927 VDPWR.n215 VDPWR.n105 17562.4
R1928 VDPWR.n217 VDPWR.n105 17562.4
R1929 VDPWR.n326 VDPWR.n323 16027.1
R1930 VDPWR.n328 VDPWR.n323 16027.1
R1931 VDPWR.n326 VDPWR.n324 16027.1
R1932 VDPWR.n328 VDPWR.n324 16027.1
R1933 VDPWR.n92 VDPWR.n89 16027.1
R1934 VDPWR.n94 VDPWR.n89 16027.1
R1935 VDPWR.n92 VDPWR.n90 16027.1
R1936 VDPWR.n94 VDPWR.n90 16027.1
R1937 VDPWR.n158 VDPWR.n142 12420
R1938 VDPWR.n158 VDPWR.n131 12420
R1939 VDPWR.n160 VDPWR.n142 12416.5
R1940 VDPWR.n160 VDPWR.n131 12416.5
R1941 VDPWR.n206 VDPWR.n119 6349.41
R1942 VDPWR.n206 VDPWR.n120 6349.41
R1943 VDPWR.n204 VDPWR.n119 6349.41
R1944 VDPWR.n204 VDPWR.n120 6349.41
R1945 VDPWR.n146 VDPWR.n141 4698.77
R1946 VDPWR.n255 VDPWR.n254 3045.88
R1947 VDPWR.n252 VDPWR.n250 3045.88
R1948 VDPWR.n254 VDPWR.n252 3045.88
R1949 VDPWR.n33 VDPWR.n30 3045.88
R1950 VDPWR.n36 VDPWR.n30 3045.88
R1951 VDPWR.n36 VDPWR.n31 3045.88
R1952 VDPWR.n310 VDPWR.n301 2701.93
R1953 VDPWR.n74 VDPWR.n9 2701.93
R1954 VDPWR.n307 VDPWR.n302 2375
R1955 VDPWR.n70 VDPWR.n11 2372.5
R1956 VDPWR.n307 VDPWR.n304 2327.31
R1957 VDPWR.n11 VDPWR.n10 2327.31
R1958 VDPWR.n279 VDPWR.n265 2089.41
R1959 VDPWR.n282 VDPWR.n264 2089.41
R1960 VDPWR.n271 VDPWR.n269 2089.41
R1961 VDPWR.n274 VDPWR.n268 2089.41
R1962 VDPWR.n286 VDPWR.n261 2089.41
R1963 VDPWR.n288 VDPWR.n246 2089.41
R1964 VDPWR.n42 VDPWR.n27 2089.41
R1965 VDPWR.n45 VDPWR.n26 2089.41
R1966 VDPWR.n49 VDPWR.n18 2089.41
R1967 VDPWR.n52 VDPWR.n17 2089.41
R1968 VDPWR.n59 VDPWR.n58 2089.41
R1969 VDPWR.n61 VDPWR.n14 2089.41
R1970 VDPWR.n179 VDPWR.n139 2071.76
R1971 VDPWR.n173 VDPWR.n164 2071.76
R1972 VDPWR.n171 VDPWR.n140 1443.53
R1973 VDPWR.n171 VDPWR.n166 1443.53
R1974 VDPWR.n328 VDPWR.t31 1353.8
R1975 VDPWR.n94 VDPWR.t19 1353.8
R1976 VDPWR.t34 VDPWR.n326 1317.74
R1977 VDPWR.t22 VDPWR.n92 1317.74
R1978 VDPWR.n327 VDPWR.t34 1196.03
R1979 VDPWR.n93 VDPWR.t22 1196.03
R1980 VDPWR.t31 VDPWR.n327 1159.97
R1981 VDPWR.t19 VDPWR.n93 1159.97
R1982 VDPWR.n167 VDPWR.n166 628.236
R1983 VDPWR.n166 VDPWR.n139 628.236
R1984 VDPWR.n173 VDPWR.n140 628.236
R1985 VDPWR.n177 VDPWR.n140 628.236
R1986 VDPWR.n237 VDPWR.n236 599.49
R1987 VDPWR.n5 VDPWR.n4 599.49
R1988 VDPWR.n325 VDPWR.n322 415.628
R1989 VDPWR.n91 VDPWR.n88 415.628
R1990 VDPWR.n72 VDPWR.t53 413.37
R1991 VDPWR.t0 VDPWR.t27 412.942
R1992 VDPWR.t17 VDPWR.t29 412.942
R1993 VDPWR.n329 VDPWR.n322 405.284
R1994 VDPWR.n95 VDPWR.n88 405.284
R1995 VDPWR.t53 VDPWR.t59 387.817
R1996 VDPWR.t27 VDPWR.n142 319.411
R1997 VDPWR.t29 VDPWR.n131 315.507
R1998 VDPWR.n280 VDPWR.n264 290.354
R1999 VDPWR.n281 VDPWR.n265 290.354
R2000 VDPWR.n272 VDPWR.n268 290.354
R2001 VDPWR.n273 VDPWR.n269 290.354
R2002 VDPWR.n288 VDPWR.n287 290.354
R2003 VDPWR.n261 VDPWR.n260 290.354
R2004 VDPWR.n43 VDPWR.n26 290.354
R2005 VDPWR.n44 VDPWR.n27 290.354
R2006 VDPWR.n50 VDPWR.n17 290.354
R2007 VDPWR.n51 VDPWR.n18 290.354
R2008 VDPWR.n61 VDPWR.n60 290.354
R2009 VDPWR.n58 VDPWR.n57 290.354
R2010 VDPWR.n305 VDPWR.n238 285.92
R2011 VDPWR.n67 VDPWR.n66 285.889
R2012 VDPWR.n71 VDPWR.n9 268.555
R2013 VDPWR.n191 VDPWR.n190 259.036
R2014 VDPWR.n306 VDPWR.n300 253.333
R2015 VDPWR.n69 VDPWR.n68 253.067
R2016 VDPWR.n309 VDPWR.n302 248.76
R2017 VDPWR.n306 VDPWR.n305 248.246
R2018 VDPWR.n68 VDPWR.n67 248.246
R2019 VDPWR.n243 VDPWR.t65 231.379
R2020 VDPWR.n20 VDPWR.t63 231.379
R2021 VDPWR.n241 VDPWR.t7 231.287
R2022 VDPWR.n293 VDPWR.t3 231.287
R2023 VDPWR.n294 VDPWR.t9 231.287
R2024 VDPWR.n81 VDPWR.t62 231.287
R2025 VDPWR.n0 VDPWR.t56 231.287
R2026 VDPWR.n22 VDPWR.t58 231.287
R2027 VDPWR.n242 VDPWR.t70 231.273
R2028 VDPWR.n21 VDPWR.t52 231.273
R2029 VDPWR.t68 VDPWR.t44 216.05
R2030 VDPWR.t13 VDPWR.t25 216.05
R2031 VDPWR.n214 VDPWR.n101 209.422
R2032 VDPWR.n159 VDPWR.t17 208.423
R2033 VDPWR.n159 VDPWR.t0 204.519
R2034 VDPWR.n295 VDPWR.n240 202.453
R2035 VDPWR.n80 VDPWR.n1 202.453
R2036 VDPWR.n325 VDPWR.n321 183.016
R2037 VDPWR.n91 VDPWR.n87 183.016
R2038 VDPWR.n303 VDPWR.n301 182.214
R2039 VDPWR.n74 VDPWR.n73 182.202
R2040 VDPWR.n254 VDPWR.t64 178.327
R2041 VDPWR.n36 VDPWR.t51 178.327
R2042 VDPWR.n330 VDPWR.n329 176.572
R2043 VDPWR.n96 VDPWR.n95 176.572
R2044 VDPWR.t11 VDPWR.n172 176.514
R2045 VDPWR.n172 VDPWR.t4 176.514
R2046 VDPWR.t44 VDPWR.n119 174.992
R2047 VDPWR.t25 VDPWR.n120 174.992
R2048 VDPWR.n250 VDPWR.n249 174.803
R2049 VDPWR.n34 VDPWR.n33 174.803
R2050 VDPWR.n179 VDPWR.n178 173.517
R2051 VDPWR.n165 VDPWR.n164 173.517
R2052 VDPWR.t15 VDPWR.n307 172.579
R2053 VDPWR.n11 VDPWR.t48 172.579
R2054 VDPWR.n175 VDPWR.n174 166.4
R2055 VDPWR.n162 VDPWR.n161 161.126
R2056 VDPWR.n219 VDPWR.n102 157.375
R2057 VDPWR.n170 VDPWR.n169 153.976
R2058 VDPWR.n170 VDPWR.n137 146.825
R2059 VDPWR.n251 VDPWR.n248 128.709
R2060 VDPWR.n37 VDPWR.n29 128.709
R2061 VDPWR.n256 VDPWR.n248 127.835
R2062 VDPWR.n168 VDPWR.n163 124.802
R2063 VDPWR.n320 VDPWR.n318 120.891
R2064 VDPWR.n86 VDPWR.n84 120.891
R2065 VDPWR.n320 VDPWR.n319 119.76
R2066 VDPWR.n86 VDPWR.n85 119.76
R2067 VDPWR.n69 VDPWR.n65 118.385
R2068 VDPWR.n311 VDPWR.n300 118.118
R2069 VDPWR.n115 VDPWR.n114 116.722
R2070 VDPWR.n218 VDPWR.n103 115.912
R2071 VDPWR.n38 VDPWR.n37 115.841
R2072 VDPWR.n219 VDPWR.n218 108.909
R2073 VDPWR.n205 VDPWR.t68 108.025
R2074 VDPWR.n205 VDPWR.t13 108.025
R2075 VDPWR.n191 VDPWR.n132 104.57
R2076 VDPWR.n270 VDPWR.n266 101.912
R2077 VDPWR.n56 VDPWR.n12 101.912
R2078 VDPWR.n136 VDPWR.t12 98.0045
R2079 VDPWR.n136 VDPWR.t5 97.6911
R2080 VDPWR.n180 VDPWR.n138 95.9841
R2081 VDPWR.n110 VDPWR.n109 87.9664
R2082 VDPWR.n110 VDPWR.n103 87.7954
R2083 VDPWR.n184 VDPWR.n135 87.2408
R2084 VDPWR.n187 VDPWR.n186 87.2408
R2085 VDPWR.n129 VDPWR.n128 87.1446
R2086 VDPWR.n151 VDPWR.n145 87.1446
R2087 VDPWR.n162 VDPWR.n141 85.5143
R2088 VDPWR.n276 VDPWR.n266 82.438
R2089 VDPWR.n56 VDPWR.n55 82.438
R2090 VDPWR.n284 VDPWR.n262 73.7015
R2091 VDPWR.n47 VDPWR.n15 73.7015
R2092 VDPWR.n277 VDPWR.n262 72.4513
R2093 VDPWR.n54 VDPWR.n15 72.4513
R2094 VDPWR.n123 VDPWR.n122 71.8902
R2095 VDPWR.t38 VDPWR.n215 71.3347
R2096 VDPWR.n203 VDPWR.n121 70.7824
R2097 VDPWR.n169 VDPWR.n168 67.0123
R2098 VDPWR.n169 VDPWR.n138 67.0123
R2099 VDPWR.n174 VDPWR.n163 65.892
R2100 VDPWR.n210 VDPWR.n106 65.6211
R2101 VDPWR.n259 VDPWR.n244 64.6513
R2102 VDPWR.n46 VDPWR.n19 64.6513
R2103 VDPWR.n259 VDPWR.n258 64.1322
R2104 VDPWR.n39 VDPWR.n19 64.1322
R2105 VDPWR.n305 VDPWR.n304 61.6672
R2106 VDPWR.n67 VDPWR.n10 61.6672
R2107 VDPWR.n174 VDPWR.n173 61.6672
R2108 VDPWR.n173 VDPWR.t11 61.6672
R2109 VDPWR.n139 VDPWR.n138 61.6672
R2110 VDPWR.t4 VDPWR.n139 61.6672
R2111 VDPWR.n168 VDPWR.n167 61.6672
R2112 VDPWR.n177 VDPWR.n176 61.6672
R2113 VDPWR.n217 VDPWR.t37 60.8049
R2114 VDPWR.n312 VDPWR.n311 58.4912
R2115 VDPWR.n65 VDPWR.n64 58.2536
R2116 VDPWR.n148 VDPWR.n147 57.394
R2117 VDPWR.n236 VDPWR.t16 57.1305
R2118 VDPWR.n236 VDPWR.t66 57.1305
R2119 VDPWR.n4 VDPWR.t49 57.1305
R2120 VDPWR.n4 VDPWR.t50 57.1305
R2121 VDPWR.n304 VDPWR.n303 56.2356
R2122 VDPWR.n73 VDPWR.n10 56.2313
R2123 VDPWR.n214 VDPWR.n213 55.3321
R2124 VDPWR.n178 VDPWR.n177 54.8697
R2125 VDPWR.n167 VDPWR.n165 54.8697
R2126 VDPWR.t43 VDPWR.t38 53.6285
R2127 VDPWR.t37 VDPWR.t10 53.6285
R2128 VDPWR.n251 VDPWR.n247 51.6747
R2129 VDPWR.n270 VDPWR.n267 51.1283
R2130 VDPWR.n207 VDPWR.n118 50.9389
R2131 VDPWR.n302 VDPWR.n300 46.2505
R2132 VDPWR.n70 VDPWR.n69 46.2505
R2133 VDPWR.n32 VDPWR.n29 45.8455
R2134 VDPWR.n308 VDPWR.t15 43.4751
R2135 VDPWR.n72 VDPWR.t48 43.4751
R2136 VDPWR.n257 VDPWR.n247 38.3351
R2137 VDPWR.n63 VDPWR.n12 36.2672
R2138 VDPWR.n157 VDPWR.n143 35.1478
R2139 VDPWR.n71 VDPWR.n70 33.6572
R2140 VDPWR.n126 VDPWR.n124 32.1789
R2141 VDPWR.t10 VDPWR.n216 32.0794
R2142 VDPWR.n126 VDPWR.n125 32.0774
R2143 VDPWR.n311 VDPWR.n310 30.8338
R2144 VDPWR.n271 VDPWR.n270 30.8338
R2145 VDPWR.n279 VDPWR.n278 30.8338
R2146 VDPWR.n275 VDPWR.n274 30.8338
R2147 VDPWR.n252 VDPWR.n251 30.8338
R2148 VDPWR.n253 VDPWR.n252 30.8338
R2149 VDPWR.n256 VDPWR.n255 30.8338
R2150 VDPWR.n246 VDPWR.n245 30.8338
R2151 VDPWR.n286 VDPWR.n285 30.8338
R2152 VDPWR.n283 VDPWR.n282 30.8338
R2153 VDPWR.n30 VDPWR.n29 30.8338
R2154 VDPWR.n35 VDPWR.n30 30.8338
R2155 VDPWR.n42 VDPWR.n41 30.8338
R2156 VDPWR.n31 VDPWR.n28 30.8338
R2157 VDPWR.n14 VDPWR.n12 30.8338
R2158 VDPWR.n65 VDPWR.n9 30.8338
R2159 VDPWR.n59 VDPWR.n13 30.8338
R2160 VDPWR.n53 VDPWR.n52 30.8338
R2161 VDPWR.n49 VDPWR.n48 30.8338
R2162 VDPWR.n46 VDPWR.n45 30.8338
R2163 VDPWR.n115 VDPWR.n106 30.7043
R2164 VDPWR.n208 VDPWR.n207 30.0503
R2165 VDPWR.n208 VDPWR.n117 29.6052
R2166 VDPWR.t59 VDPWR.n71 29.2303
R2167 VDPWR.n255 VDPWR.n249 28.7736
R2168 VDPWR.n34 VDPWR.n31 28.7736
R2169 VDPWR.n240 VDPWR.t42 28.5655
R2170 VDPWR.n240 VDPWR.t40 28.5655
R2171 VDPWR.n1 VDPWR.t60 28.5655
R2172 VDPWR.n1 VDPWR.t54 28.5655
R2173 VDPWR.n280 VDPWR.n279 26.1635
R2174 VDPWR.n272 VDPWR.n271 26.1635
R2175 VDPWR.n274 VDPWR.n273 26.1635
R2176 VDPWR.n287 VDPWR.n286 26.1635
R2177 VDPWR.n260 VDPWR.n246 26.1635
R2178 VDPWR.n282 VDPWR.n281 26.1635
R2179 VDPWR.n43 VDPWR.n42 26.1635
R2180 VDPWR.n50 VDPWR.n49 26.1635
R2181 VDPWR.n52 VDPWR.n51 26.1635
R2182 VDPWR.n60 VDPWR.n59 26.1635
R2183 VDPWR.n57 VDPWR.n14 26.1635
R2184 VDPWR.n45 VDPWR.n44 26.1635
R2185 VDPWR.n148 VDPWR.n146 24.2792
R2186 VDPWR.n310 VDPWR.n309 23.2602
R2187 VDPWR.n268 VDPWR.n266 23.1311
R2188 VDPWR.n58 VDPWR.n56 23.1311
R2189 VDPWR.n264 VDPWR.n262 23.1255
R2190 VDPWR.n269 VDPWR.n267 23.1255
R2191 VDPWR.n265 VDPWR.n263 23.1255
R2192 VDPWR.n261 VDPWR.n259 23.1255
R2193 VDPWR.n289 VDPWR.n288 23.1255
R2194 VDPWR.n26 VDPWR.n19 23.1255
R2195 VDPWR.n40 VDPWR.n27 23.1255
R2196 VDPWR.n18 VDPWR.n15 23.1255
R2197 VDPWR.n62 VDPWR.n61 23.1255
R2198 VDPWR.n17 VDPWR.n16 23.1255
R2199 VDPWR.n41 VDPWR.n40 22.5272
R2200 VDPWR.n216 VDPWR.t43 21.5497
R2201 VDPWR.n164 VDPWR.n163 18.5005
R2202 VDPWR.n180 VDPWR.n179 18.5005
R2203 VDPWR.n171 VDPWR.n170 18.5005
R2204 VDPWR.n172 VDPWR.n171 18.5005
R2205 VDPWR.n32 VDPWR.n28 18.4652
R2206 VDPWR.n181 VDPWR.n180 18.1802
R2207 VDPWR.n181 VDPWR.n137 17.9947
R2208 VDPWR.n257 VDPWR.n256 16.1646
R2209 VDPWR.n319 VDPWR.t36 15.8699
R2210 VDPWR.n319 VDPWR.t32 15.8699
R2211 VDPWR.n318 VDPWR.t35 15.8699
R2212 VDPWR.n318 VDPWR.t33 15.8699
R2213 VDPWR.n85 VDPWR.t24 15.8699
R2214 VDPWR.n85 VDPWR.t21 15.8699
R2215 VDPWR.n84 VDPWR.t23 15.8699
R2216 VDPWR.n84 VDPWR.t20 15.8699
R2217 VDPWR.n313 VDPWR.n312 14.6418
R2218 VDPWR.n76 VDPWR.n3 14.6377
R2219 VDPWR.n298 VDPWR.n238 14.5701
R2220 VDPWR.n66 VDPWR.n8 14.5701
R2221 VDPWR.n283 VDPWR.n263 12.9491
R2222 VDPWR.n275 VDPWR.n267 12.7742
R2223 VDPWR.n278 VDPWR.n263 12.7334
R2224 VDPWR.n313 VDPWR.n299 12.7275
R2225 VDPWR.n76 VDPWR.n75 12.7273
R2226 VDPWR.n289 VDPWR.n245 12.6169
R2227 VDPWR.n290 VDPWR.n289 12.3941
R2228 VDPWR.n64 VDPWR.n63 12.0598
R2229 VDPWR.n161 VDPWR.n133 11.6663
R2230 VDPWR.n307 VDPWR.n306 11.563
R2231 VDPWR.n68 VDPWR.n11 11.563
R2232 VDPWR.n135 VDPWR.t28 11.4265
R2233 VDPWR.n135 VDPWR.t47 11.4265
R2234 VDPWR.n186 VDPWR.t18 11.4265
R2235 VDPWR.n186 VDPWR.t30 11.4265
R2236 VDPWR.n128 VDPWR.t67 11.4265
R2237 VDPWR.n128 VDPWR.t46 11.4265
R2238 VDPWR.n145 VDPWR.t41 11.4265
R2239 VDPWR.n145 VDPWR.t1 11.4265
R2240 VDPWR.n277 VDPWR.n276 11.3214
R2241 VDPWR.n285 VDPWR.n284 11.0119
R2242 VDPWR.n254 VDPWR.n248 10.8829
R2243 VDPWR.n250 VDPWR.n247 10.8829
R2244 VDPWR.n37 VDPWR.n36 10.8829
R2245 VDPWR.n33 VDPWR.n32 10.8829
R2246 VDPWR.n63 VDPWR.n62 10.3636
R2247 VDPWR.n329 VDPWR.n328 10.2783
R2248 VDPWR.n326 VDPWR.n325 10.2783
R2249 VDPWR.n95 VDPWR.n94 10.2783
R2250 VDPWR.n92 VDPWR.n91 10.2783
R2251 VDPWR.n48 VDPWR.n16 9.97982
R2252 VDPWR.n62 VDPWR.n13 9.86377
R2253 VDPWR.n55 VDPWR.n54 9.85683
R2254 VDPWR.n53 VDPWR.n16 9.83647
R2255 VDPWR.n73 VDPWR.n72 9.79085
R2256 VDPWR.n308 VDPWR.n303 9.78762
R2257 VDPWR.n39 VDPWR.n38 9.73877
R2258 VDPWR.n312 VDPWR.n239 9.68315
R2259 VDPWR.n78 VDPWR.n3 9.6823
R2260 VDPWR.n47 VDPWR.n46 9.62493
R2261 VDPWR.n40 VDPWR.n25 9.59483
R2262 VDPWR.n6 VDPWR 9.58101
R2263 VDPWR.n114 VDPWR.n113 9.34567
R2264 VDPWR.n144 VDPWR.n143 9.3005
R2265 VDPWR.n154 VDPWR.n132 9.3005
R2266 VDPWR.n134 VDPWR.n133 9.3005
R2267 VDPWR.n202 VDPWR.n201 9.3005
R2268 VDPWR.n211 VDPWR.n210 9.3005
R2269 VDPWR.n111 VDPWR.n110 9.3005
R2270 VDPWR.n309 VDPWR.t39 9.2139
R2271 VDPWR.n258 VDPWR.n257 9.03689
R2272 VDPWR.t64 VDPWR.n253 8.9954
R2273 VDPWR.t51 VDPWR.n35 8.9954
R2274 VDPWR.n122 VDPWR.n120 8.04398
R2275 VDPWR.n121 VDPWR.n119 8.04398
R2276 VDPWR.n301 VDPWR.n299 7.4005
R2277 VDPWR.n75 VDPWR.n74 7.4005
R2278 VDPWR.n295 VDPWR 7.28043
R2279 VDPWR VDPWR.n80 7.20708
R2280 VDPWR.n204 VDPWR.n203 7.11588
R2281 VDPWR.n205 VDPWR.n204 7.11588
R2282 VDPWR.n207 VDPWR.n206 7.11588
R2283 VDPWR.n206 VDPWR.n205 7.11588
R2284 VDPWR.n213 VDPWR.n106 6.56253
R2285 VDPWR.n176 VDPWR.n175 5.75273
R2286 VDPWR.n192 VDPWR.n131 5.60656
R2287 VDPWR.n147 VDPWR.n142 5.60656
R2288 VDPWR.n109 VDPWR.n105 5.44168
R2289 VDPWR.n216 VDPWR.n105 5.44168
R2290 VDPWR.n104 VDPWR.n102 5.44168
R2291 VDPWR.n216 VDPWR.n104 5.44168
R2292 VDPWR.t11 VDPWR.n165 5.16575
R2293 VDPWR.n178 VDPWR.t4 5.16575
R2294 VDPWR.n317 VDPWR 4.92656
R2295 VDPWR.n203 VDPWR.n202 4.82369
R2296 VDPWR.n175 VDPWR.n162 4.58844
R2297 VDPWR.t39 VDPWR.n308 4.5733
R2298 VDPWR.n154 VDPWR.n153 4.5005
R2299 VDPWR.n185 VDPWR.n134 4.5005
R2300 VDPWR.n121 VDPWR.n118 4.48345
R2301 VDPWR.n114 VDPWR.n107 4.42232
R2302 VDPWR.n281 VDPWR.t2 4.28573
R2303 VDPWR.n273 VDPWR.t8 4.28573
R2304 VDPWR.t8 VDPWR.n272 4.28573
R2305 VDPWR.t2 VDPWR.n280 4.28573
R2306 VDPWR.n260 VDPWR.t6 4.28573
R2307 VDPWR.n287 VDPWR.t6 4.28573
R2308 VDPWR.n44 VDPWR.t57 4.28573
R2309 VDPWR.t57 VDPWR.n43 4.28573
R2310 VDPWR.n57 VDPWR.t61 4.28573
R2311 VDPWR.n60 VDPWR.t61 4.28573
R2312 VDPWR.n51 VDPWR.t55 4.28573
R2313 VDPWR.t55 VDPWR.n50 4.28573
R2314 VDPWR.n124 VDPWR.t45 4.08121
R2315 VDPWR.n124 VDPWR.t69 4.08121
R2316 VDPWR.n125 VDPWR.t14 4.08121
R2317 VDPWR.n125 VDPWR.t26 4.08121
R2318 VDPWR.n196 VDPWR.n127 3.98496
R2319 VDPWR.n189 VDPWR.n130 3.8313
R2320 VDPWR.n227 VDPWR 3.4738
R2321 VDPWR.n228 VDPWR 3.41826
R2322 VDPWR.n147 VDPWR.n141 3.22115
R2323 VDPWR.n229 VDPWR 3.19356
R2324 VDPWR.n182 VDPWR.n134 3.09113
R2325 VDPWR.n161 VDPWR.n160 2.68166
R2326 VDPWR.n160 VDPWR.n159 2.68166
R2327 VDPWR.n158 VDPWR.n157 2.68166
R2328 VDPWR.n159 VDPWR.n158 2.68166
R2329 VDPWR.n187 VDPWR.n127 2.55635
R2330 VDPWR.n232 VDPWR 2.21561
R2331 VDPWR.n83 VDPWR 2.1638
R2332 VDPWR.n234 VDPWR 2.12067
R2333 VDPWR.n202 VDPWR.n123 1.94833
R2334 VDPWR.n235 VDPWR.n82 1.91485
R2335 VDPWR.n113 VDPWR.n112 1.87667
R2336 VDPWR.n109 VDPWR.n107 1.86232
R2337 VDPWR.n195 VDPWR.n194 1.85463
R2338 VDPWR.n222 VDPWR.n221 1.85361
R2339 VDPWR.n154 VDPWR.n130 1.78294
R2340 VDPWR.n253 VDPWR.n249 1.7705
R2341 VDPWR.n35 VDPWR.n34 1.7705
R2342 VDPWR.n333 VDPWR.n332 1.75798
R2343 VDPWR.n184 VDPWR.n183 1.688
R2344 VDPWR.n215 VDPWR.n214 1.66717
R2345 VDPWR.n218 VDPWR.n217 1.66717
R2346 VDPWR.n324 VDPWR.n322 1.63767
R2347 VDPWR.n327 VDPWR.n324 1.63767
R2348 VDPWR.n323 VDPWR.n321 1.63767
R2349 VDPWR.n327 VDPWR.n323 1.63767
R2350 VDPWR.n90 VDPWR.n88 1.63767
R2351 VDPWR.n93 VDPWR.n90 1.63767
R2352 VDPWR.n89 VDPWR.n87 1.63767
R2353 VDPWR.n93 VDPWR.n89 1.63767
R2354 VDPWR.n24 VDPWR.n20 1.62503
R2355 VDPWR.n291 VDPWR.n243 1.6242
R2356 VDPWR.n209 VDPWR.n208 1.6211
R2357 VDPWR.n190 VDPWR.n133 1.45873
R2358 VDPWR.n185 VDPWR.n184 1.27935
R2359 VDPWR.n331 VDPWR 1.27612
R2360 VDPWR.n97 VDPWR 1.27612
R2361 VDPWR.n99 VDPWR.n98 1.23754
R2362 VDPWR.n317 VDPWR 1.22297
R2363 VDPWR.n102 VDPWR.n101 1.20392
R2364 VDPWR.n332 VDPWR.n320 1.20189
R2365 VDPWR.n98 VDPWR.n86 1.20189
R2366 VDPWR.n122 VDPWR.n117 1.19816
R2367 VDPWR.n149 VDPWR.n144 1.19668
R2368 VDPWR.n156 VDPWR.n132 1.19015
R2369 VDPWR.n334 VDPWR 1.17597
R2370 VDPWR.n149 VDPWR.n148 1.11733
R2371 VDPWR.n231 VDPWR 1.05905
R2372 VDPWR.n146 VDPWR.n143 1.05462
R2373 VDPWR.n234 VDPWR.n233 1.04215
R2374 VDPWR.n294 VDPWR.n293 1.01465
R2375 VDPWR.n242 VDPWR.n241 1.00136
R2376 VDPWR.n22 VDPWR.n21 1.00136
R2377 VDPWR.n212 VDPWR.n211 0.985286
R2378 VDPWR.n224 VDPWR.n99 0.96796
R2379 VDPWR.n111 VDPWR.n108 0.96321
R2380 VDPWR.n188 VDPWR.n187 0.963107
R2381 VDPWR.n176 VDPWR.n137 0.933293
R2382 VDPWR.n200 VDPWR.n199 0.928261
R2383 VDPWR.n233 VDPWR.n232 0.913357
R2384 VDPWR.n212 VDPWR.n115 0.875256
R2385 VDPWR.n213 VDPWR.n212 0.862026
R2386 VDPWR.n220 VDPWR.n100 0.84882
R2387 VDPWR.n197 VDPWR.n196 0.838031
R2388 VDPWR.n317 VDPWR.n235 0.833105
R2389 VDPWR.n77 VDPWR.n7 0.813514
R2390 VDPWR.n315 VDPWR.n314 0.813496
R2391 VDPWR.n155 VDPWR.n144 0.780009
R2392 VDPWR.n112 VDPWR.n111 0.758322
R2393 VDPWR.n299 VDPWR.n298 0.649348
R2394 VDPWR.n75 VDPWR.n8 0.649348
R2395 VDPWR.n150 VDPWR.n149 0.641762
R2396 VDPWR.n223 VDPWR.n100 0.634469
R2397 VDPWR.n23 VDPWR.n22 0.612135
R2398 VDPWR.n292 VDPWR.n241 0.611349
R2399 VDPWR.n192 VDPWR.n191 0.603552
R2400 VDPWR.n292 VDPWR.n291 0.595437
R2401 VDPWR.n24 VDPWR.n23 0.595437
R2402 VDPWR.n182 VDPWR.n181 0.58175
R2403 VDPWR.n198 VDPWR.n197 0.539263
R2404 VDPWR.n82 VDPWR.n0 0.529588
R2405 VDPWR.n330 VDPWR.n321 0.492808
R2406 VDPWR.n96 VDPWR.n87 0.492808
R2407 VDPWR.n230 VDPWR 0.464203
R2408 VDPWR.n199 VDPWR.n198 0.445398
R2409 VDPWR.n233 VDPWR 0.430018
R2410 VDPWR.n195 VDPWR.n129 0.41511
R2411 VDPWR.n151 VDPWR.n150 0.407233
R2412 VDPWR.n293 VDPWR.n292 0.403802
R2413 VDPWR.n23 VDPWR.n0 0.403016
R2414 VDPWR.n314 VDPWR.n313 0.358192
R2415 VDPWR.n77 VDPWR.n76 0.358192
R2416 VDPWR.n152 VDPWR.n151 0.347903
R2417 VDPWR.n112 VDPWR.n103 0.342518
R2418 VDPWR.n315 VDPWR.n238 0.332643
R2419 VDPWR.n66 VDPWR.n7 0.332643
R2420 VDPWR.n197 VDPWR.n118 0.321789
R2421 VDPWR.n243 VDPWR.n242 0.319213
R2422 VDPWR.n21 VDPWR.n20 0.319213
R2423 VDPWR.n153 VDPWR.n129 0.314461
R2424 VDPWR.n235 VDPWR 0.282694
R2425 VDPWR.n227 VDPWR.n226 0.263348
R2426 VDPWR.n157 VDPWR.n156 0.2565
R2427 VDPWR.n183 VDPWR.n182 0.2505
R2428 VDPWR.n284 VDPWR.n283 0.242713
R2429 VDPWR.n298 VDPWR.n297 0.239152
R2430 VDPWR.n8 VDPWR.n2 0.239152
R2431 VDPWR.n64 VDPWR.n3 0.237537
R2432 VDPWR.n229 VDPWR.n228 0.233738
R2433 VDPWR.n38 VDPWR.n28 0.228778
R2434 VDPWR.n224 VDPWR.n223 0.224984
R2435 VDPWR.n48 VDPWR.n47 0.212205
R2436 VDPWR VDPWR.n316 0.182446
R2437 VDPWR.n82 VDPWR.n81 0.180531
R2438 VDPWR.n220 VDPWR.n99 0.167373
R2439 VDPWR.n225 VDPWR.n224 0.164719
R2440 VDPWR.n79 VDPWR.n2 0.163235
R2441 VDPWR.n297 VDPWR.n296 0.162905
R2442 VDPWR.n296 VDPWR.n239 0.1505
R2443 VDPWR.n316 VDPWR.n315 0.1505
R2444 VDPWR.n79 VDPWR.n78 0.1505
R2445 VDPWR.n7 VDPWR.n6 0.1505
R2446 VDPWR.n193 VDPWR.n192 0.1505
R2447 VDPWR.n190 VDPWR.n189 0.148119
R2448 VDPWR.n210 VDPWR.n209 0.137839
R2449 VDPWR.n183 VDPWR.n136 0.133423
R2450 VDPWR.n290 VDPWR.n244 0.130922
R2451 VDPWR.n108 VDPWR.n107 0.129667
R2452 VDPWR.n199 VDPWR.n117 0.129667
R2453 VDPWR.n331 VDPWR.n330 0.123496
R2454 VDPWR.n97 VDPWR.n96 0.123496
R2455 VDPWR.n46 VDPWR.n25 0.114495
R2456 VDPWR.n297 VDPWR.n237 0.112307
R2457 VDPWR.n5 VDPWR.n2 0.111978
R2458 VDPWR.n200 VDPWR.n123 0.103833
R2459 VDPWR.n221 VDPWR.n219 0.0994362
R2460 VDPWR.n258 VDPWR.n245 0.0936587
R2461 VDPWR.n226 VDPWR 0.0868949
R2462 VDPWR.n222 VDPWR.n101 0.0866111
R2463 VDPWR.n54 VDPWR.n53 0.0831873
R2464 VDPWR.n41 VDPWR.n39 0.0819249
R2465 VDPWR VDPWR.n334 0.0802064
R2466 VDPWR.n278 VDPWR.n277 0.0763519
R2467 VDPWR.n291 VDPWR.n290 0.0678913
R2468 VDPWR.n25 VDPWR.n24 0.0678913
R2469 VDPWR.n194 VDPWR.n193 0.0666765
R2470 VDPWR.n189 VDPWR.n188 0.0638803
R2471 VDPWR.n232 VDPWR.n83 0.0578659
R2472 VDPWR.n276 VDPWR.n275 0.0573889
R2473 VDPWR VDPWR.n294 0.0571038
R2474 VDPWR.n81 VDPWR 0.0571038
R2475 VDPWR.n221 VDPWR.n220 0.0566005
R2476 VDPWR.n6 VDPWR.n5 0.0519512
R2477 VDPWR.n316 VDPWR.n237 0.0516214
R2478 VDPWR.n55 VDPWR.n13 0.0501124
R2479 VDPWR.n228 VDPWR.n227 0.0473828
R2480 VDPWR.n201 VDPWR.n126 0.047375
R2481 VDPWR.n150 VDPWR 0.0443375
R2482 VDPWR.n234 VDPWR.n83 0.0382175
R2483 VDPWR.n223 VDPWR.n222 0.038
R2484 VDPWR.n78 VDPWR.n77 0.037915
R2485 VDPWR.n314 VDPWR.n239 0.0370646
R2486 VDPWR.n196 VDPWR.n195 0.0364015
R2487 VDPWR.n209 VDPWR.n116 0.0341957
R2488 VDPWR.n296 VDPWR.n295 0.0303556
R2489 VDPWR.n80 VDPWR.n79 0.0303556
R2490 VDPWR.n156 VDPWR.n155 0.0274565
R2491 VDPWR.n155 VDPWR.n154 0.0266936
R2492 VDPWR.n153 VDPWR.n152 0.0261494
R2493 VDPWR.n194 VDPWR.n127 0.0233659
R2494 VDPWR.n201 VDPWR.n200 0.0216694
R2495 VDPWR.n189 VDPWR.n134 0.0211422
R2496 VDPWR.n198 VDPWR.n116 0.020648
R2497 VDPWR.n188 VDPWR.n185 0.0197308
R2498 VDPWR.n285 VDPWR.n244 0.0191317
R2499 VDPWR.n193 VDPWR.n130 0.0144018
R2500 VDPWR.n332 VDPWR.n331 0.0133125
R2501 VDPWR.n98 VDPWR.n97 0.0133125
R2502 VDPWR.n155 VDPWR.n152 0.0121883
R2503 VDPWR.n235 VDPWR.n234 0.00943855
R2504 VDPWR.n233 VDPWR.n231 0.00624391
R2505 VDPWR.n231 VDPWR.n230 0.00363011
R2506 VDPWR.n211 VDPWR.n116 0.00255592
R2507 VDPWR.n333 VDPWR.n317 0.00209349
R2508 VDPWR.n334 VDPWR.n333 0.00209349
R2509 VDPWR.n113 VDPWR.n108 0.00155302
R2510 VDPWR.n226 VDPWR.n225 0.00104613
R2511 VDPWR.n100 VDPWR 0.000994071
R2512 VDPWR.n225 VDPWR 0.000663025
R2513 VDPWR.n230 VDPWR.n229 0.000568264
R2514 a_24889_22946.t0 a_24889_22946.t1 50.1091
R2515 3_OTA_0.OTA_stage1_0.vd1 3_OTA_0.OTA_stage1_0.vd1.t2 122.216
R2516 3_OTA_0.OTA_stage1_0.vd1 3_OTA_0.OTA_stage1_0.vd1.t3 122.216
R2517 3_OTA_0.OTA_stage1_0.vd1 3_OTA_0.OTA_stage1_0.vd1.t0 121.828
R2518 3_OTA_0.OTA_stage1_0.vd1 3_OTA_0.OTA_stage1_0.vd1.t1 121.828
R2519 a_3013_4521.t19 a_3013_4521.n39 190.305
R2520 a_3013_4521.n43 a_3013_4521.t19 190.305
R2521 a_3013_4521.t33 a_3013_4521.n41 190.305
R2522 a_3013_4521.n42 a_3013_4521.t33 190.305
R2523 a_3013_4521.n34 a_3013_4521.t29 190.305
R2524 a_3013_4521.t29 a_3013_4521.n24 190.305
R2525 a_3013_4521.t39 a_3013_4521.n35 190.305
R2526 a_3013_4521.n36 a_3013_4521.t39 190.305
R2527 a_3013_4521.t31 a_3013_4521.n47 190.305
R2528 a_3013_4521.n51 a_3013_4521.t31 190.305
R2529 a_3013_4521.t37 a_3013_4521.n49 190.305
R2530 a_3013_4521.n50 a_3013_4521.t37 190.305
R2531 a_3013_4521.t15 a_3013_4521.n17 190.305
R2532 a_3013_4521.n12 a_3013_4521.t15 190.305
R2533 a_3013_4521.t21 a_3013_4521.n62 190.305
R2534 a_3013_4521.n63 a_3013_4521.t21 190.305
R2535 a_3013_4521.n58 a_3013_4521.t27 190.305
R2536 a_3013_4521.n20 a_3013_4521.t27 190.305
R2537 a_3013_4521.t41 a_3013_4521.n19 190.305
R2538 a_3013_4521.n55 a_3013_4521.t41 190.305
R2539 a_3013_4521.t23 a_3013_4521.n71 190.305
R2540 a_3013_4521.n72 a_3013_4521.t23 190.305
R2541 a_3013_4521.t13 a_3013_4521.n69 190.305
R2542 a_3013_4521.n73 a_3013_4521.t13 190.305
R2543 a_3013_4521.t25 a_3013_4521.n80 190.305
R2544 a_3013_4521.n81 a_3013_4521.t25 190.305
R2545 a_3013_4521.t43 a_3013_4521.n14 190.305
R2546 a_3013_4521.n82 a_3013_4521.t43 190.305
R2547 a_3013_4521.n78 a_3013_4521.t35 95.1811
R2548 a_3013_4521.n23 a_3013_4521.t17 95.1783
R2549 a_3013_4521.n22 a_3013_4521.n21 22.3176
R2550 a_3013_4521.n67 a_3013_4521.n66 22.2301
R2551 a_3013_4521.n27 a_3013_4521.n26 22.2284
R2552 a_3013_4521.n9 a_3013_4521.n28 22.2284
R2553 a_3013_4521.n31 a_3013_4521.n30 22.2284
R2554 a_3013_4521.n11 a_3013_4521.n29 22.2284
R2555 a_3013_4521.n5 a_3013_4521.n68 22.2284
R2556 a_3013_4521.n0 a_3013_4521.n75 22.2284
R2557 a_3013_4521.n7 a_3013_4521.n76 22.2284
R2558 a_3013_4521.n6 a_3013_4521.n45 22.1884
R2559 a_3013_4521.n10 a_3013_4521.n46 22.1884
R2560 a_3013_4521.n2 a_3013_4521.n53 22.1884
R2561 a_3013_4521.n3 a_3013_4521.n54 22.1884
R2562 a_3013_4521.n1 a_3013_4521.n13 22.1884
R2563 a_3013_4521.n4 a_3013_4521.n77 22.1884
R2564 a_3013_4521.n84 a_3013_4521.n8 22.1884
R2565 a_3013_4521.n38 a_3013_4521.n23 11.5981
R2566 a_3013_4521.n79 a_3013_4521.n78 10.9335
R2567 a_3013_4521.n80 a_3013_4521.n79 9.89233
R2568 a_3013_4521.n39 a_3013_4521.n38 9.80925
R2569 a_3013_4521.n47 a_3013_4521.n18 9.80925
R2570 a_3013_4521.n59 a_3013_4521.n58 9.80925
R2571 a_3013_4521.n73 a_3013_4521.n16 9.48127
R2572 a_3013_4521.n12 a_3013_4521.n60 9.40378
R2573 a_3013_4521.n37 a_3013_4521.n36 9.39819
R2574 a_3013_4521.n27 a_3013_4521.n23 4.9275
R2575 a_3013_4521.n78 a_3013_4521.n7 4.79654
R2576 a_3013_4521.n0 a_3013_4521.n74 4.5005
R2577 a_3013_4521.n70 a_3013_4521.n5 4.5005
R2578 a_3013_4521.n65 a_3013_4521.n64 4.5005
R2579 a_3013_4521.n61 a_3013_4521.n11 4.5005
R2580 a_3013_4521.n32 a_3013_4521.n25 4.5005
R2581 a_3013_4521.n33 a_3013_4521.n9 4.5005
R2582 a_3013_4521.n15 a_3013_4521.n4 4.5005
R2583 a_3013_4521.n8 a_3013_4521.n83 4.5005
R2584 a_3013_4521.n3 a_3013_4521.n56 4.5005
R2585 a_3013_4521.n57 a_3013_4521.n1 4.5005
R2586 a_3013_4521.n48 a_3013_4521.n10 4.5005
R2587 a_3013_4521.n2 a_3013_4521.n52 4.5005
R2588 a_3013_4521.n40 a_3013_4521.n22 4.5005
R2589 a_3013_4521.n6 a_3013_4521.n44 4.5005
R2590 a_3013_4521.n21 a_3013_4521.t7 4.3505
R2591 a_3013_4521.n21 a_3013_4521.t34 4.3505
R2592 a_3013_4521.n45 a_3013_4521.t20 4.3505
R2593 a_3013_4521.n45 a_3013_4521.t4 4.3505
R2594 a_3013_4521.n46 a_3013_4521.t1 4.3505
R2595 a_3013_4521.n46 a_3013_4521.t38 4.3505
R2596 a_3013_4521.n53 a_3013_4521.t32 4.3505
R2597 a_3013_4521.n53 a_3013_4521.t45 4.3505
R2598 a_3013_4521.n54 a_3013_4521.t3 4.3505
R2599 a_3013_4521.n54 a_3013_4521.t42 4.3505
R2600 a_3013_4521.n13 a_3013_4521.t28 4.3505
R2601 a_3013_4521.n13 a_3013_4521.t0 4.3505
R2602 a_3013_4521.n77 a_3013_4521.t26 4.3505
R2603 a_3013_4521.n77 a_3013_4521.t8 4.3505
R2604 a_3013_4521.n26 a_3013_4521.t18 4.3505
R2605 a_3013_4521.n26 a_3013_4521.t47 4.3505
R2606 a_3013_4521.n28 a_3013_4521.t10 4.3505
R2607 a_3013_4521.n28 a_3013_4521.t30 4.3505
R2608 a_3013_4521.n30 a_3013_4521.t40 4.3505
R2609 a_3013_4521.n30 a_3013_4521.t2 4.3505
R2610 a_3013_4521.n29 a_3013_4521.t12 4.3505
R2611 a_3013_4521.n29 a_3013_4521.t22 4.3505
R2612 a_3013_4521.n66 a_3013_4521.t16 4.3505
R2613 a_3013_4521.n66 a_3013_4521.t5 4.3505
R2614 a_3013_4521.n68 a_3013_4521.t11 4.3505
R2615 a_3013_4521.n68 a_3013_4521.t24 4.3505
R2616 a_3013_4521.n75 a_3013_4521.t14 4.3505
R2617 a_3013_4521.n75 a_3013_4521.t46 4.3505
R2618 a_3013_4521.n76 a_3013_4521.t6 4.3505
R2619 a_3013_4521.n76 a_3013_4521.t36 4.3505
R2620 a_3013_4521.n84 a_3013_4521.t9 4.3505
R2621 a_3013_4521.t44 a_3013_4521.n84 4.3505
R2622 a_3013_4521.n7 a_3013_4521.n4 2.55258
R2623 a_3013_4521.n38 a_3013_4521.n37 1.86108
R2624 a_3013_4521.n37 a_3013_4521.n18 1.86108
R2625 a_3013_4521.n60 a_3013_4521.n18 1.86108
R2626 a_3013_4521.n60 a_3013_4521.n59 1.86108
R2627 a_3013_4521.n59 a_3013_4521.n16 1.86108
R2628 a_3013_4521.n79 a_3013_4521.n16 1.86108
R2629 a_3013_4521.n7 a_3013_4521.n0 1.20675
R2630 a_3013_4521.n9 a_3013_4521.n27 1.0755
R2631 a_3013_4521.n31 a_3013_4521.n11 1.0755
R2632 a_3013_4521.n5 a_3013_4521.n67 1.0755
R2633 a_3013_4521.n10 a_3013_4521.n6 1.0755
R2634 a_3013_4521.n3 a_3013_4521.n2 1.0755
R2635 a_3013_4521.n8 a_3013_4521.n1 1.0755
R2636 a_3013_4521.n62 a_3013_4521.n61 0.759759
R2637 a_3013_4521.n64 a_3013_4521.n17 0.756673
R2638 a_3013_4521.n35 a_3013_4521.n25 0.702205
R2639 a_3013_4521.n34 a_3013_4521.n33 0.700784
R2640 a_3013_4521.n56 a_3013_4521.n55 0.669534
R2641 a_3013_4521.n52 a_3013_4521.n51 0.668114
R2642 a_3013_4521.n44 a_3013_4521.n43 0.666693
R2643 a_3013_4521.n57 a_3013_4521.n20 0.665273
R2644 a_3013_4521.n83 a_3013_4521.n82 0.662432
R2645 a_3013_4521.n81 a_3013_4521.n15 0.661011
R2646 a_3013_4521.n42 a_3013_4521.n40 0.659208
R2647 a_3013_4521.n64 a_3013_4521.n12 0.647608
R2648 a_3013_4521.n63 a_3013_4521.n61 0.645562
R2649 a_3013_4521.n80 a_3013_4521.n15 0.632599
R2650 a_3013_4521.n83 a_3013_4521.n14 0.631182
R2651 a_3013_4521.n50 a_3013_4521.n48 0.629532
R2652 a_3013_4521.n58 a_3013_4521.n57 0.628338
R2653 a_3013_4521.n44 a_3013_4521.n39 0.626917
R2654 a_3013_4521.n52 a_3013_4521.n47 0.625497
R2655 a_3013_4521.n56 a_3013_4521.n19 0.62408
R2656 a_3013_4521.n41 a_3013_4521.n40 0.619882
R2657 a_3013_4521.n49 a_3013_4521.n48 0.594586
R2658 a_3013_4521.n33 a_3013_4521.n24 0.59283
R2659 a_3013_4521.n36 a_3013_4521.n25 0.591408
R2660 a_3013_4521.n74 a_3013_4521.n69 0.580689
R2661 a_3013_4521.n71 a_3013_4521.n70 0.57833
R2662 a_3013_4521.n2 a_3013_4521.n10 0.538
R2663 a_3013_4521.n1 a_3013_4521.n3 0.538
R2664 a_3013_4521.n0 a_3013_4521.n5 0.538
R2665 a_3013_4521.n8 a_3013_4521.n4 0.536231
R2666 a_3013_4521.n72 a_3013_4521.n70 0.495783
R2667 a_3013_4521.n74 a_3013_4521.n73 0.493424
R2668 a_3013_4521.n12 a_3013_4521.n63 0.488952
R2669 a_3013_4521.n62 a_3013_4521.n17 0.486913
R2670 a_3013_4521.n41 a_3013_4521.n39 0.476043
R2671 a_3013_4521.n43 a_3013_4521.n42 0.476043
R2672 a_3013_4521.n49 a_3013_4521.n47 0.459739
R2673 a_3013_4521.n51 a_3013_4521.n50 0.459739
R2674 a_3013_4521.n58 a_3013_4521.n19 0.459739
R2675 a_3013_4521.n55 a_3013_4521.n20 0.459739
R2676 a_3013_4521.n80 a_3013_4521.n14 0.459739
R2677 a_3013_4521.n82 a_3013_4521.n81 0.459739
R2678 a_3013_4521.n36 a_3013_4521.n24 0.451587
R2679 a_3013_4521.n35 a_3013_4521.n34 0.451587
R2680 a_3013_4521.n6 a_3013_4521.n22 0.408833
R2681 a_3013_4521.n73 a_3013_4521.n72 0.405391
R2682 a_3013_4521.n71 a_3013_4521.n69 0.405391
R2683 a_3013_4521.n65 a_3013_4521.n11 0.395292
R2684 a_3013_4521.n9 a_3013_4521.n32 0.395292
R2685 a_3013_4521.n32 a_3013_4521.n31 0.143208
R2686 a_3013_4521.n67 a_3013_4521.n65 0.143208
R2687 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 936.04
R2688 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 235.982
R2689 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 235.978
R2690 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 190.305
R2691 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 190.305
R2692 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 190.305
R2693 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 190.305
R2694 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 190.305
R2695 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 190.305
R2696 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 95.3928
R2697 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 95.3656
R2698 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 95.1789
R2699 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 95.1648
R2700 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 95.1535
R2701 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 95.1535
R2702 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 94.8314
R2703 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 94.8314
R2704 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 94.8314
R2705 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 94.8314
R2706 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 94.8314
R2707 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 94.8314
R2708 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 94.8314
R2709 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 94.8314
R2710 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 94.8314
R2711 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 94.8314
R2712 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 94.8314
R2713 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 94.8314
R2714 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 94.8314
R2715 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 94.8314
R2716 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 94.8314
R2717 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 94.8314
R2718 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 94.8314
R2719 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 94.8314
R2720 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 94.8314
R2721 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 94.8314
R2722 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 94.8314
R2723 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 94.8314
R2724 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 94.8314
R2725 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 84.0884
R2726 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 83.5719
R2727 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 83.5719
R2728 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 83.5719
R2729 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 83.5719
R2730 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 73.19
R2731 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 26.074
R2732 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 26.074
R2733 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 26.074
R2734 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 25.7843
R2735 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 10.2824
R2736 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 9.66398
R2737 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R2738 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R2739 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R2740 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R2741 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R2742 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R2743 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R2744 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R2745 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R2746 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R2747 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R2748 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R2749 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R2750 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R2751 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R2752 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 9.3005
R2753 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 9.3005
R2754 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R2755 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 9.3005
R2756 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R2757 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R2758 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R2759 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R2760 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R2761 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 9.3005
R2762 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R2763 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R2764 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 9.3005
R2765 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 7.22993
R2766 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 7.22993
R2767 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 7.20169
R2768 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 6.83022
R2769 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 6.81633
R2770 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 6.81633
R2771 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 6.81633
R2772 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 6.75312
R2773 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 4.64588
R2774 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 4.64588
R2775 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 4.64588
R2776 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 4.64588
R2777 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 2.29815
R2778 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 1.86108
R2779 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 1.86108
R2780 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 1.86108
R2781 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 1.86108
R2782 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 1.86108
R2783 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 1.86108
R2784 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 1.86108
R2785 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 1.28691
R2786 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 1.25468
R2787 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 1.14402
R2788 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 1.1424
R2789 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 1.12066
R2790 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 1.12066
R2791 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 1.11251
R2792 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 1.10979
R2793 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 1.10164
R2794 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 1.10164
R2795 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 1.10164
R2796 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 1.10164
R2797 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 1.09892
R2798 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 1.09349
R2799 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 1.09349
R2800 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 1.08805
R2801 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 1.08262
R2802 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 1.08262
R2803 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 1.08262
R2804 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 1.07024
R2805 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 1.0237
R2806 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.959578
R2807 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 0.812055
R2808 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.77514
R2809 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.701365
R2810 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.645119
R2811 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 0.645119
R2812 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 0.645119
R2813 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 0.645119
R2814 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 0.645119
R2815 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 0.645119
R2816 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 0.645119
R2817 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.645119
R2818 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 0.645119
R2819 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.645119
R2820 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 0.645119
R2821 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 0.645119
R2822 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 0.645119
R2823 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 0.645119
R2824 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 0.645119
R2825 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.645119
R2826 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 0.645119
R2827 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.645119
R2828 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 0.645119
R2829 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 0.645119
R2830 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 0.645119
R2831 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 0.645119
R2832 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 0.645119
R2833 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.645119
R2834 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.645119
R2835 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 0.645119
R2836 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 0.645119
R2837 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 0.645119
R2838 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 0.645119
R2839 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 0.645118
R2840 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 0.590702
R2841 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 0.572258
R2842 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 0.495065
R2843 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.495065
R2844 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 0.481478
R2845 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.481478
R2846 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.475521
R2847 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 0.470609
R2848 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.470609
R2849 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 0.465174
R2850 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 0.465174
R2851 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.465174
R2852 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.459844
R2853 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 0.459739
R2854 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.459739
R2855 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 0.446152
R2856 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.446152
R2857 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.445943
R2858 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.443435
R2859 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.440717
R2860 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 0.440717
R2861 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.434551
R2862 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 0.432313
R2863 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.414484
R2864 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.408265
R2865 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.408265
R2866 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.40372
R2867 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.40372
R2868 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.314045
R2869 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 0.290206
R2870 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 0.0183279
R2871 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 0.0112346
R2872 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 0.0112346
R2873 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.0112346
R2874 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 0.0112346
R2875 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.0112346
R2876 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 0.0112346
R2877 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 0.0112346
R2878 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 0.0112346
R2879 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 0.00760547
R2880 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 0.00316393
R2881 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t0 88.7532
R2882 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n14 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n12 22.2005
R2883 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n3 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n1 21.8665
R2884 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n26 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n25 21.5445
R2885 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n24 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n23 21.5445
R2886 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n22 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n21 21.5445
R2887 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n20 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n19 21.5445
R2888 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n18 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n17 21.5445
R2889 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n16 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n15 21.5445
R2890 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n14 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n13 21.5445
R2891 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n11 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n10 21.5445
R2892 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n9 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n8 21.5445
R2893 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n7 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n6 21.5445
R2894 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n5 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n4 21.5445
R2895 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n3 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n2 21.5445
R2896 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n0 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n29 21.5445
R2897 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n28 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n27 21.5418
R2898 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n27 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t22 4.3505
R2899 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n27 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t11 4.3505
R2900 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n25 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t32 4.3505
R2901 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n25 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t25 4.3505
R2902 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n23 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t20 4.3505
R2903 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n23 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t12 4.3505
R2904 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n21 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t31 4.3505
R2905 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n21 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t15 4.3505
R2906 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n19 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t19 4.3505
R2907 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n19 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t10 4.3505
R2908 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n17 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t2 4.3505
R2909 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n17 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t16 4.3505
R2910 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n15 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t18 4.3505
R2911 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n15 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t5 4.3505
R2912 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n13 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t30 4.3505
R2913 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n13 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t21 4.3505
R2914 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n12 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t17 4.3505
R2915 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n12 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t13 4.3505
R2916 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n10 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t23 4.3505
R2917 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n10 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t9 4.3505
R2918 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n8 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t6 4.3505
R2919 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n8 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t28 4.3505
R2920 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n6 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t24 4.3505
R2921 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n6 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t1 4.3505
R2922 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n4 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t3 4.3505
R2923 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n4 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t27 4.3505
R2924 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n2 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t14 4.3505
R2925 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n2 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t8 4.3505
R2926 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n1 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t4 4.3505
R2927 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n1 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t26 4.3505
R2928 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n29 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t7 4.3505
R2929 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n29 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t29 4.3505
R2930 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n28 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n26 1.51316
R2931 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n18 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n16 0.624699
R2932 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n22 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n20 0.624699
R2933 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n26 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n24 0.624699
R2934 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n5 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n3 0.60872
R2935 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n9 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n7 0.60872
R2936 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n0 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n11 0.553215
R2937 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n0 0.408658
R2938 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n0 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n28 0.298079
R2939 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n16 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n14 0.296969
R2940 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n20 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n18 0.296969
R2941 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n24 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n22 0.296969
R2942 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n7 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n5 0.289615
R2943 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n11 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n9 0.289615
R2944 3_OTA_0.OTA_vref_0.vb1.n1 3_OTA_0.OTA_vref_0.vb1.n2 71.7516
R2945 3_OTA_0.OTA_vref_0.vb1.n1 3_OTA_0.OTA_vref_0.vb1.n4 70.9453
R2946 3_OTA_0.OTA_vref_0.vb1.n1 3_OTA_0.OTA_vref_0.vb1.n3 70.9453
R2947 3_OTA_0.OTA_vref_0.vb1.n0 3_OTA_0.OTA_vref_0.vb1.t9 68.1062
R2948 3_OTA_0.OTA_vref_0.vb1.n0 3_OTA_0.OTA_vref_0.vb1.t7 67.5138
R2949 3_OTA_0.OTA_vref_0.vb1.n0 3_OTA_0.OTA_vref_0.vb1.t8 67.5138
R2950 3_OTA_0.OTA_vref_0.vb1.n0 3_OTA_0.OTA_vref_0.vb1.t6 67.5138
R2951 3_OTA_0.OTA_vref_0.vb1.n2 3_OTA_0.OTA_vref_0.vb1.t0 17.4005
R2952 3_OTA_0.OTA_vref_0.vb1.n2 3_OTA_0.OTA_vref_0.vb1.t3 17.4005
R2953 3_OTA_0.OTA_vref_0.vb1.n4 3_OTA_0.OTA_vref_0.vb1.t2 17.4005
R2954 3_OTA_0.OTA_vref_0.vb1.n4 3_OTA_0.OTA_vref_0.vb1.t1 17.4005
R2955 3_OTA_0.OTA_vref_0.vb1.n3 3_OTA_0.OTA_vref_0.vb1.t5 17.4005
R2956 3_OTA_0.OTA_vref_0.vb1.n3 3_OTA_0.OTA_vref_0.vb1.t4 17.4005
R2957 3_OTA_0.OTA_vref_0.vb1 3_OTA_0.OTA_vref_0.vb1.n0 10.0205
R2958 3_OTA_0.OTA_vref_0.vb1 3_OTA_0.OTA_vref_0.vb1.n1 8.74264
R2959 a_12564_25551.n8 a_12564_25551.t11 36.4777
R2960 a_12564_25551.n7 a_12564_25551.t8 35.4327
R2961 a_12564_25551.n9 a_12564_25551.n8 31.3519
R2962 a_12564_25551.n5 a_12564_25551.n4 18.3035
R2963 a_12564_25551.n2 a_12564_25551.n1 18.303
R2964 a_12564_25551.n5 a_12564_25551.n3 17.2098
R2965 a_12564_25551.n2 a_12564_25551.n0 17.208
R2966 a_12564_25551.n6 a_12564_25551.n2 8.938
R2967 a_12564_25551.n9 a_12564_25551.t9 4.08121
R2968 a_12564_25551.t10 a_12564_25551.n9 4.08121
R2969 a_12564_25551.n6 a_12564_25551.n5 3.05142
R2970 a_12564_25551.n7 a_12564_25551.n6 2.2455
R2971 a_12564_25551.n4 a_12564_25551.t3 1.90483
R2972 a_12564_25551.n4 a_12564_25551.t7 1.90483
R2973 a_12564_25551.n3 a_12564_25551.t0 1.90483
R2974 a_12564_25551.n3 a_12564_25551.t4 1.90483
R2975 a_12564_25551.n1 a_12564_25551.t6 1.90483
R2976 a_12564_25551.n1 a_12564_25551.t5 1.90483
R2977 a_12564_25551.n0 a_12564_25551.t2 1.90483
R2978 a_12564_25551.n0 a_12564_25551.t1 1.90483
R2979 a_12564_25551.n8 a_12564_25551.n7 1.0455
R2980 3_OTA_0.3rd_3_OTA_0.vd4.n2 3_OTA_0.3rd_3_OTA_0.vd4.t10 82.3324
R2981 3_OTA_0.3rd_3_OTA_0.vd4.n0 3_OTA_0.3rd_3_OTA_0.vd4.t11 81.6762
R2982 3_OTA_0.3rd_3_OTA_0.vd4.n2 3_OTA_0.3rd_3_OTA_0.vd4.t12 81.6762
R2983 3_OTA_0.3rd_3_OTA_0.vd4.n0 3_OTA_0.3rd_3_OTA_0.vd4.t8 81.4249
R2984 3_OTA_0.3rd_3_OTA_0.vd4.n6 3_OTA_0.3rd_3_OTA_0.vd4.t4 72.7606
R2985 3_OTA_0.3rd_3_OTA_0.vd4.n1 3_OTA_0.3rd_3_OTA_0.vd4.t5 71.6732
R2986 3_OTA_0.3rd_3_OTA_0.vd4 3_OTA_0.3rd_3_OTA_0.vd4.n7 62.243
R2987 3_OTA_0.3rd_3_OTA_0.vd4.n4 3_OTA_0.3rd_3_OTA_0.vd4.t3 19.4751
R2988 3_OTA_0.3rd_3_OTA_0.vd4.n4 3_OTA_0.3rd_3_OTA_0.vd4.t2 18.6511
R2989 3_OTA_0.3rd_3_OTA_0.vd4.n5 3_OTA_0.3rd_3_OTA_0.vd4.n3 15.6099
R2990 3_OTA_0.3rd_3_OTA_0.vd4.n7 3_OTA_0.3rd_3_OTA_0.vd4.t7 11.6005
R2991 3_OTA_0.3rd_3_OTA_0.vd4.n7 3_OTA_0.3rd_3_OTA_0.vd4.t6 11.6005
R2992 3_OTA_0.3rd_3_OTA_0.vd4.n1 3_OTA_0.3rd_3_OTA_0.vd4.t9 4.23179
R2993 3_OTA_0.3rd_3_OTA_0.vd4.n1 3_OTA_0.3rd_3_OTA_0.vd4.n6 2.48505
R2994 3_OTA_0.3rd_3_OTA_0.vd4.n3 3_OTA_0.3rd_3_OTA_0.vd4.t0 1.90483
R2995 3_OTA_0.3rd_3_OTA_0.vd4.n3 3_OTA_0.3rd_3_OTA_0.vd4.t1 1.90483
R2996 3_OTA_0.3rd_3_OTA_0.vd4 3_OTA_0.3rd_3_OTA_0.vd4.n0 1.4105
R2997 3_OTA_0.3rd_3_OTA_0.vd4.n5 3_OTA_0.3rd_3_OTA_0.vd4.n4 1.32214
R2998 3_OTA_0.3rd_3_OTA_0.vd4.n6 3_OTA_0.3rd_3_OTA_0.vd4.n5 1.28407
R2999 3_OTA_0.3rd_3_OTA_0.vd4.n0 3_OTA_0.3rd_3_OTA_0.vd4.n2 0.8105
R3000 3_OTA_0.3rd_3_OTA_0.vd4 3_OTA_0.3rd_3_OTA_0.vd4.n1 0.42303
R3001 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd2.t3 134.761
R3002 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd2.t2 134.73
R3003 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd2.t4 122.688
R3004 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd2.t5 122.213
R3005 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd2.t6 122.213
R3006 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd2.t7 121.831
R3007 3_OTA_0.OTA_stage1_0.vd2.t0 3_OTA_0.OTA_stage1_0.vd2.t1 27.306
R3008 ua[1].n0 ua[1].t0 138.714
R3009 ua[1].n2 ua[1].t1 136.073
R3010 ua[1].n0 ua[1].t2 19.5045
R3011 ua[1].n1 ua[1].t3 17.559
R3012 ua[1].n1 ua[1].n0 6.3305
R3013 ua[1].n2 ua[1].n1 1.803
R3014 ua[1] ua[1].n2 0.337827
R3015 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n0 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t17 651.943
R3016 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n18 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t19 651.74
R3017 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n20 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t24 60.1752
R3018 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n19 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t22 60.1752
R3019 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n10 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t0 28.5589
R3020 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n14 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t10 27.6016
R3021 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n21 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t23 26.8562
R3022 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n21 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t26 26.0492
R3023 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n22 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t21 26.0492
R3024 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n23 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t25 26.0492
R3025 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n24 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t20 26.0492
R3026 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n5 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n4 24.2089
R3027 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n11 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n8 23.2516
R3028 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n10 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n9 23.2516
R3029 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n7 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n1 23.2516
R3030 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n6 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n2 23.2516
R3031 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n5 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n3 23.2516
R3032 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n13 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n12 23.2516
R3033 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n17 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t18 23
R3034 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n0 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t16 23
R3035 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n8 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t13 4.3505
R3036 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n8 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t9 4.3505
R3037 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n9 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t14 4.3505
R3038 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n9 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t7 4.3505
R3039 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n1 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t6 4.3505
R3040 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n1 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t1 4.3505
R3041 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n2 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t8 4.3505
R3042 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n2 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t5 4.3505
R3043 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n3 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t11 4.3505
R3044 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n3 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t4 4.3505
R3045 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n4 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t12 4.3505
R3046 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n4 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t3 4.3505
R3047 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n12 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t15 4.3505
R3048 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n12 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t2 4.3505
R3049 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n16 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n15 3.8934
R3050 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n22 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n21 2.80213
R3051 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n24 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n23 2.76952
R3052 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n23 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n22 2.72333
R3053 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n15 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n7 1.06728
R3054 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n7 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n6 0.957816
R3055 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n6 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n5 0.957816
R3056 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n14 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n13 0.957816
R3057 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n13 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n11 0.957816
R3058 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n11 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n10 0.957816
R3059 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n19 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n18 0.712457
R3060 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n20 0.660826
R3061 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n24 0.617348
R3062 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n15 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n14 0.577487
R3063 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n20 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n19 0.36463
R3064 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n17 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n16 0.240192
R3065 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n16 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n0 0.216951
R3066 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n18 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n17 0.206939
R3067 ua[0].n0 ua[0].t0 98.4603
R3068 ua[0].n0 ua[0].t2 88.6727
R3069 ua[0].n1 ua[0].t1 46.53
R3070 ua[0].n1 ua[0].n0 0.203972
R3071 ua[0] ua[0].n1 0.107444
R3072 ua[3].n1 ua[3].t0 21.0692
R3073 ua[3].n0 ua[3].t1 21.0692
R3074 ua[3] ua[3].n2 10.0582
R3075 ua[3].n1 ua[3].t3 8.85313
R3076 ua[3].n0 ua[3].t2 8.85313
R3077 ua[3] ua[3].n1 2.40005
R3078 ua[3] ua[3].n0 2.40005
R3079 ua[3].n2 ua[3] 1.67184
R3080 ua[3].n2 ua[3] 0.685917
R3081 a_21048_25880.n8 a_21048_25880.t12 387.724
R3082 a_21048_25880.n7 a_21048_25880.t9 96.3265
R3083 a_21048_25880.n4 a_21048_25880.t5 96.3265
R3084 a_21048_25880.n0 a_21048_25880.n9 84.9005
R3085 a_21048_25880.n3 a_21048_25880.t2 38.5275
R3086 a_21048_25880.t3 a_21048_25880.n3 37.908
R3087 a_21048_25880.n3 a_21048_25880.n10 32.1023
R3088 a_21048_25880.n4 a_21048_25880.n5 0.971171
R3089 a_21048_25880.n7 a_21048_25880.n6 0.710684
R3090 a_21048_25880.n0 a_21048_25880.t6 13.2778
R3091 a_21048_25880.n1 a_21048_25880.n0 1.6868
R3092 a_21048_25880.n6 a_21048_25880.t8 13.6521
R3093 a_21048_25880.n1 a_21048_25880.t10 12.8838
R3094 a_21048_25880.t4 a_21048_25880.n5 13.4238
R3095 a_21048_25880.n9 a_21048_25880.t11 11.4265
R3096 a_21048_25880.n9 a_21048_25880.t7 11.4265
R3097 a_21048_25880.n0 a_21048_25880.n3 6.81377
R3098 a_21048_25880.n3 a_21048_25880.n4 6.43072
R3099 a_21048_25880.n2 a_21048_25880.n1 4.23945
R3100 a_21048_25880.n10 a_21048_25880.t0 5.8005
R3101 a_21048_25880.n10 a_21048_25880.t1 5.8005
R3102 a_21048_25880.n8 a_21048_25880.n2 0.713738
R3103 a_21048_25880.n2 a_21048_25880.n6 9.2977
R3104 a_21048_25880.n5 a_21048_25880.n8 6.84764
R3105 a_21048_25880.n7 a_21048_25880.n3 6.18407
R3106 a_21048_27042.n9 a_21048_27042.t12 387.31
R3107 a_21048_27042.n10 a_21048_27042.t11 96.3265
R3108 a_21048_27042.n6 a_21048_27042.t7 96.3265
R3109 a_21048_27042.n3 a_21048_27042.n8 84.9005
R3110 a_21048_27042.t3 a_21048_27042.n5 35.0885
R3111 a_21048_27042.n5 a_21048_27042.t2 34.5018
R3112 a_21048_27042.t10 a_21048_27042.n9 32.649
R3113 a_21048_27042.n7 a_21048_27042.n6 0.971171
R3114 a_21048_27042.n10 a_21048_27042.t10 28.9361
R3115 a_21048_27042.n5 a_21048_27042.n11 28.9216
R3116 a_21048_27042.t8 a_21048_27042.n3 28.1453
R3117 a_21048_27042.n2 a_21048_27042.t4 13.2766
R3118 a_21048_27042.n7 a_21048_27042.t6 13.4238
R3119 a_21048_27042.n8 a_21048_27042.t5 11.4265
R3120 a_21048_27042.n8 a_21048_27042.t9 11.4265
R3121 a_21048_27042.n0 a_21048_27042.n7 7.07514
R3122 a_21048_27042.n1 a_21048_27042.n0 2.67922
R3123 a_21048_27042.n11 a_21048_27042.t0 5.8005
R3124 a_21048_27042.n11 a_21048_27042.t1 5.8005
R3125 a_21048_27042.n1 a_21048_27042.n2 1.64285
R3126 a_21048_27042.n4 a_21048_27042.n6 5.19734
R3127 a_21048_27042.n5 a_21048_27042.n3 3.73846
R3128 a_21048_27042.n9 a_21048_27042.n0 3.7305
R3129 a_21048_27042.n4 a_21048_27042.n10 3.46037
R3130 a_21048_27042.n2 a_21048_27042.n3 1.08359
R3131 a_21048_27042.n5 a_21048_27042.n4 1.8052
R3132 a_21048_27042.n1 a_21048_27042.t8 27.348
R3133 ua[5].n4 ua[5].t5 231.043
R3134 ua[5].n3 ua[5].t3 85.987
R3135 ua[5].n2 ua[5].n0 71.7516
R3136 ua[5].n2 ua[5].n1 70.9453
R3137 ua[5].n0 ua[5].t4 17.4005
R3138 ua[5].n0 ua[5].t2 17.4005
R3139 ua[5].n1 ua[5].t1 17.4005
R3140 ua[5].n1 ua[5].t0 17.4005
R3141 ua[5].n3 ua[5].n2 0.896828
R3142 ua[5].n4 ua[5].n3 0.859275
R3143 ua[5] ua[5].n4 0.129667
R3144 ua[4] ua[4].t0 15.4738
C0 3_OTA_0.OTA_vref_0.vb a_22654_21988# 0.541253f
C1 ua[2] 3_OTA_0.OTA_vref_0.vb 0.408082f
C2 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter VDPWR 0.504763f
C3 a_16084_17427# a_15996_17227# 1.53765f
C4 a_15996_21097# VDPWR 0.368035f
C5 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 a_15996_17227# 0.112341f
C6 3_OTA_0.3rd_3_OTA_0.vd3 a_15996_21097# 0.001347f
C7 3_OTA_0.OTA_stage1_0.vd1 a_25461_23684# 0.011993f
C8 a_15996_21097# 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.002329f
C9 ua[4] a_18046_7223# 0.440838f
C10 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 2.20693f
C11 VDPWR a_16084_17427# 0.034292f
C12 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 VDPWR 0.030224f
C13 a_6631_3101# a_6631_4391# 0.154422f
C14 a_16084_17427# 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.003419f
C15 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 16.2573f
C16 3_OTA_0.3rd_3_OTA_0.vd4 3_OTA_0.OTA_vref_0.vb1 0.226739f
C17 VDPWR a_16084_20007# 0.034455f
C18 a_6631_6971# BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 0.112195f
C19 ua[3] VDPWR 0.335831f
C20 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_16084_20007# 6.62e-20
C21 ua[3] a_18046_7223# 1.47482f
C22 a_6631_4391# BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 0.334532f
C23 a_6719_6913# BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.002793f
C24 3_OTA_0.OTA_vref_0.vb a_3537_27009# 0.443825f
C25 a_15996_17227# a_15996_18517# 0.154705f
C26 3_OTA_0.OTA_stage1_0.vd1 VDPWR 8.443541f
C27 a_6719_4333# VDPWR 0.034455f
C28 a_6719_5623# BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 1.65e-19
C29 3_OTA_0.3rd_3_OTA_0.vd4 a_15996_21097# 2.1e-20
C30 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.OTA_stage1_0.vd1 1.22886f
C31 ua[2] a_3537_27009# 1.68092f
C32 VDPWR a_15996_18517# 0.318981f
C33 a_6631_5681# BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 0.011611f
C34 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_15996_18517# 0.009524f
C35 a_6631_5681# a_6631_4391# 0.154516f
C36 ua[5] ua[3] 0.076108f
C37 VDPWR a_25461_23684# 0.836592f
C38 3_OTA_0.3rd_3_OTA_0.vd3 a_25461_23684# 6.67e-20
C39 3_OTA_0.3rd_3_OTA_0.vd4 3_OTA_0.OTA_stage1_0.vd1 15.7657f
C40 a_6719_5623# a_6719_4333# 0.036353f
C41 ua[2] ua[1] 0.138779f
C42 ua[5] a_6719_4333# 0.036384f
C43 3_OTA_0.OTA_stage1_0.vd1 ua[0] 0.367637f
C44 VDPWR a_15996_17227# 0.3278f
C45 a_6631_3101# BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 0.367242f
C46 a_15996_17227# 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.032619f
C47 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 16.257f
C48 3_OTA_0.3rd_3_OTA_0.vd3 VDPWR 4.64542f
C49 3_OTA_0.OTA_vref_0.vb1 a_15996_19807# 0.106848f
C50 a_18046_7223# VDPWR 5.64e-19
C51 VDPWR 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.512021f
C52 3_OTA_0.3rd_3_OTA_0.vd4 a_25461_23684# 1.15e-20
C53 a_6631_4391# BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.005854f
C54 3_OTA_0.OTA_vref_0.vb 3_OTA_0.OTA_vref_0.vb1 0.111837f
C55 a_6631_6971# BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 0.335671f
C56 ua[0] a_25461_23684# 0.159655f
C57 a_15996_21097# a_15996_19807# 0.154422f
C58 a_6719_6913# VDPWR 0.034292f
C59 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 a_6719_4333# 0.001293f
C60 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 a_15996_19807# 0.011315f
C61 a_6719_5623# VDPWR 0.034493f
C62 3_OTA_0.3rd_3_OTA_0.vd4 VDPWR 4.41784f
C63 3_OTA_0.OTA_vref_0.vb a_15996_21097# 1.67298f
C64 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.3rd_3_OTA_0.vd4 9.480929f
C65 a_16084_20007# a_15996_19807# 1.53005f
C66 a_6631_5681# BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 0.340876f
C67 ua[5] VDPWR 0.31178f
C68 3_OTA_0.OTA_vref_0.vb 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 4.32e-19
C69 ua[0] VDPWR 3.17609f
C70 a_6631_4391# a_6719_4333# 1.53005f
C71 ua[4] ua[2] 0.328127f
C72 a_6631_6971# a_6631_5681# 0.154705f
C73 3_OTA_0.OTA_vref_0.vb a_16084_20007# 0.036384f
C74 ua[3] 3_OTA_0.OTA_vref_0.vb 0.618087f
C75 a_6719_6913# a_6719_5623# 0.036353f
C76 a_15996_19807# a_15996_18517# 0.154516f
C77 ua[2] ua[3] 5.69043f
C78 3_OTA_0.OTA_vref_0.vb 3_OTA_0.OTA_stage1_0.vd1 0.2466f
C79 a_6631_3101# BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 5.07e-19
C80 3_OTA_0.OTA_stage1_0.vd1 a_22654_21988# 0.006984f
C81 ua[2] 3_OTA_0.OTA_stage1_0.vd1 0.13787f
C82 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 9.25527f
C83 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 VDPWR 0.030808f
C84 ua[3] a_3537_27009# 1.47482f
C85 a_6631_6971# BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.024292f
C86 ua[4] ua[1] 0.200778f
C87 a_6631_4391# VDPWR 0.335621f
C88 3_OTA_0.OTA_stage1_0.vd1 a_3537_27009# 0.118468f
C89 a_22654_21988# a_25461_23684# 0.016974f
C90 a_6631_3101# a_6719_4333# 0.10061f
C91 VDPWR a_15996_19807# 0.335707f
C92 a_6719_6913# BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 0.037992f
C93 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_15996_19807# 0.007176f
C94 ua[3] ua[1] 0.784618f
C95 a_6719_4333# BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 0.008037f
C96 a_6631_5681# BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.00639f
C97 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 a_6719_5623# 0.001618f
C98 3_OTA_0.OTA_vref_0.vb VDPWR 0.434712f
C99 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.OTA_vref_0.vb 0.136282f
C100 3_OTA_0.OTA_vref_0.vb 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.006315f
C101 VDPWR a_22654_21988# 0.101608f
C102 ua[2] VDPWR 0.298348f
C103 3_OTA_0.3rd_3_OTA_0.vd3 a_22654_21988# 1.06971f
C104 a_6719_5623# a_6631_4391# 0.098772f
C105 ua[2] a_18046_7223# 1.68131f
C106 ua[5] a_6631_4391# 3.04e-19
C107 a_6631_5681# a_6719_4333# 1.04e-19
C108 3_OTA_0.OTA_vref_0.vb 3_OTA_0.3rd_3_OTA_0.vd4 0.001057f
C109 a_16084_17427# 3_OTA_0.OTA_vref_0.vb1 0.056235f
C110 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 3_OTA_0.OTA_vref_0.vb1 0.006422f
C111 a_3537_27009# VDPWR 5.64e-19
C112 3_OTA_0.OTA_vref_0.vb1 a_16084_20007# 0.038035f
C113 a_6631_3101# VDPWR 0.369319f
C114 3_OTA_0.3rd_3_OTA_0.vd4 a_22654_21988# 1.05152f
C115 VDPWR BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 11.3779f
C116 ua[0] a_22654_21988# 0.004168f
C117 a_15996_21097# a_16084_20007# 0.10061f
C118 a_6631_6971# VDPWR 0.324581f
C119 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 a_16084_17427# 0.037994f
C120 3_OTA_0.OTA_vref_0.vb1 a_15996_18517# 1.61373f
C121 ua[1] VDPWR 2.53878f
C122 ua[4] ua[3] 0.734728f
C123 a_18046_7223# ua[1] 0.118468f
C124 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 a_16084_20007# 0.00151f
C125 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 a_6631_4391# 0.01076f
C126 a_6719_4333# BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 1.58e-19
C127 a_6719_6913# BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 0.008049f
C128 ua[5] a_6631_3101# 1.6531f
C129 a_6719_5623# BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 0.008143f
C130 a_6631_6971# a_6719_6913# 1.53765f
C131 a_6631_5681# VDPWR 0.318904f
C132 a_16084_17427# a_15996_18517# 0.097592f
C133 ua[5] BGR_BJT_vref_0.BGR_BJT_stage2_0.vr 0.174409f
C134 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 a_15996_18517# 0.010991f
C135 ua[3] 3_OTA_0.OTA_stage1_0.vd1 0.784618f
C136 a_6631_6971# a_6719_5623# 1.04e-19
C137 a_16084_20007# a_15996_18517# 1.04e-19
C138 a_15996_17227# 3_OTA_0.OTA_vref_0.vb1 0.034229f
C139 3_OTA_0.OTA_vref_0.vb a_15996_19807# 3.04e-19
C140 a_6719_6913# a_6631_5681# 0.097608f
C141 VDPWR 3_OTA_0.OTA_vref_0.vb1 8.322209f
C142 3_OTA_0.3rd_3_OTA_0.vd3 3_OTA_0.OTA_vref_0.vb1 0.316815f
C143 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 3_OTA_0.OTA_vref_0.vb1 6.15e-19
C144 a_6631_5681# a_6719_5623# 1.53781f
C145 ua[4] VGND 8.86421f
C146 ua[5] VGND 3.78062f
C147 ua[1] VGND 14.056011f
C148 ua[0] VGND 16.261526f
C149 ua[3] VGND 47.99248f
C150 ua[2] VGND 47.096302f
C151 VDPWR VGND 36.89474f
C152 a_18046_7223# VGND 3.49104f
C153 a_6631_3101# VGND 3.74629f
C154 a_6719_4333# VGND 0.471213f
C155 a_6631_4391# VGND 3.71343f
C156 a_6719_5623# VGND 0.471213f
C157 a_6631_5681# VGND 3.71408f
C158 a_6719_6913# VGND 0.471596f
C159 a_6631_6971# VGND 3.84028f
C160 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0 VGND 9.207773f
C161 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter VGND 25.328465f
C162 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr VGND 12.144946f
C163 a_15996_17227# VGND 3.83372f
C164 a_16084_17427# VGND 0.471548f
C165 a_15996_18517# VGND 3.70817f
C166 a_15996_19807# VGND 3.70757f
C167 a_16084_20007# VGND 0.471213f
C168 a_15996_21097# VGND 3.74966f
C169 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0 VGND 9.084187f
C170 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter VGND 25.297863f
C171 a_25461_23684# VGND 1.4749f
C172 a_22654_21988# VGND 5.75308f
C173 3_OTA_0.OTA_vref_0.vb1 VGND 8.843204f
C174 3_OTA_0.3rd_3_OTA_0.vd3 VGND 50.17144f
C175 3_OTA_0.3rd_3_OTA_0.vd4 VGND 19.390491f
C176 3_OTA_0.OTA_vref_0.vb VGND 18.3013f
C177 a_3537_27009# VGND 3.49104f
C178 3_OTA_0.OTA_stage1_0.vd1 VGND 84.930405f
C179 a_21048_27042.n0 VGND 1.17962f
C180 a_21048_27042.n1 VGND 1.22804f
C181 a_21048_27042.n2 VGND 0.281253f
C182 a_21048_27042.t4 VGND 1.50909f
C183 a_21048_27042.n3 VGND 1.29217f
C184 a_21048_27042.n4 VGND 1.58696f
C185 a_21048_27042.n5 VGND 3.86795f
C186 a_21048_27042.n6 VGND 1.02899f
C187 a_21048_27042.n7 VGND 0.64178f
C188 a_21048_27042.t12 VGND 0.12612f
C189 a_21048_27042.t7 VGND 0.081856f
C190 a_21048_27042.t6 VGND 1.51857f
C191 a_21048_27042.t5 VGND 0.022262f
C192 a_21048_27042.t9 VGND 0.022262f
C193 a_21048_27042.n8 VGND 0.045353f
C194 a_21048_27042.t8 VGND 1.52061f
C195 a_21048_27042.n9 VGND 1.63593f
C196 a_21048_27042.t10 VGND 1.63702f
C197 a_21048_27042.t11 VGND 0.081856f
C198 a_21048_27042.n10 VGND 0.711803f
C199 a_21048_27042.t0 VGND 0.026714f
C200 a_21048_27042.t1 VGND 0.026714f
C201 a_21048_27042.n11 VGND 0.078485f
C202 a_21048_27042.t2 VGND 0.118908f
C203 a_21048_27042.t3 VGND 0.129672f
C204 a_21048_25880.n0 VGND 1.46343f
C205 a_21048_25880.n1 VGND 0.936679f
C206 a_21048_25880.n2 VGND 1.29294f
C207 a_21048_25880.n3 VGND 5.4296f
C208 a_21048_25880.n4 VGND 0.906851f
C209 a_21048_25880.n5 VGND 0.620305f
C210 a_21048_25880.n6 VGND 0.742801f
C211 a_21048_25880.n7 VGND 0.763129f
C212 a_21048_25880.n8 VGND 1.26286f
C213 a_21048_25880.t2 VGND 0.150205f
C214 a_21048_25880.t12 VGND 0.127287f
C215 a_21048_25880.t8 VGND 1.5052f
C216 a_21048_25880.t9 VGND 0.080806f
C217 a_21048_25880.t6 VGND 1.48973f
C218 a_21048_25880.t11 VGND 0.021976f
C219 a_21048_25880.t7 VGND 0.021976f
C220 a_21048_25880.n9 VGND 0.044771f
C221 a_21048_25880.t10 VGND 1.48363f
C222 a_21048_25880.t4 VGND 1.49909f
C223 a_21048_25880.t5 VGND 0.080806f
C224 a_21048_25880.t0 VGND 0.026371f
C225 a_21048_25880.t1 VGND 0.026371f
C226 a_21048_25880.n10 VGND 0.083184f
C227 a_21048_25880.t3 VGND 0.13999f
C228 ua[3].t1 VGND 0.765616f
C229 ua[3].t2 VGND 0.402811f
C230 ua[3].n0 VGND 0.887113f
C231 ua[3].t0 VGND 0.765614f
C232 ua[3].t3 VGND 0.402811f
C233 ua[3].n1 VGND 0.887116f
C234 ua[3].n2 VGND 0.736438f
C235 ua[0].t1 VGND 0.009938f
C236 ua[0].t0 VGND 0.016128f
C237 ua[0].t2 VGND 0.006215f
C238 ua[0].n0 VGND 0.070622f
C239 ua[0].n1 VGND 0.107769f
C240 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t24 VGND 0.303177f
C241 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t22 VGND 0.303177f
C242 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t19 VGND 0.025819f
C243 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t17 VGND 0.025848f
C244 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t16 VGND 0.458348f
C245 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n0 VGND 0.831668f
C246 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t6 VGND 0.054701f
C247 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t1 VGND 0.054701f
C248 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n1 VGND 0.207792f
C249 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t8 VGND 0.054701f
C250 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t5 VGND 0.054701f
C251 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n2 VGND 0.207792f
C252 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t11 VGND 0.054701f
C253 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t4 VGND 0.054701f
C254 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n3 VGND 0.207792f
C255 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t12 VGND 0.054701f
C256 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t3 VGND 0.054701f
C257 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n4 VGND 0.236001f
C258 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n5 VGND 1.66404f
C259 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n6 VGND 0.978905f
C260 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n7 VGND 1.01624f
C261 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t10 VGND 0.275825f
C262 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t13 VGND 0.054701f
C263 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t9 VGND 0.054701f
C264 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n8 VGND 0.207792f
C265 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t14 VGND 0.054701f
C266 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t7 VGND 0.054701f
C267 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n9 VGND 0.207792f
C268 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t0 VGND 0.301124f
C269 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n10 VGND 1.70832f
C270 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n11 VGND 0.978905f
C271 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t15 VGND 0.054701f
C272 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t2 VGND 0.054701f
C273 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n12 VGND 0.207792f
C274 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n13 VGND 0.978905f
C275 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n14 VGND 0.920186f
C276 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n15 VGND 1.6821f
C277 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n16 VGND 0.842958f
C278 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t18 VGND 0.458348f
C279 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n17 VGND 0.767751f
C280 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n18 VGND 0.122062f
C281 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n19 VGND 0.367555f
C282 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n20 VGND 0.365494f
C283 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t23 VGND 0.607306f
C284 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t26 VGND 0.584001f
C285 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n21 VGND 1.65121f
C286 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t21 VGND 0.584001f
C287 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n22 VGND 0.975491f
C288 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t25 VGND 0.584001f
C289 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n23 VGND 0.974189f
C290 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.t20 VGND 0.584001f
C291 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr.n24 VGND 0.890133f
C292 ua[1].t1 VGND 0.049297f
C293 ua[1].t0 VGND 0.054519f
C294 ua[1].t2 VGND 0.405248f
C295 ua[1].n0 VGND 2.2097f
C296 ua[1].t3 VGND 0.247711f
C297 ua[1].n1 VGND 1.41396f
C298 ua[1].n2 VGND 0.590676f
C299 3_OTA_0.OTA_stage1_0.vd2.t0 VGND 38.682198f
C300 3_OTA_0.OTA_stage1_0.vd2.t4 VGND 1.331f
C301 3_OTA_0.OTA_stage1_0.vd2.t6 VGND 1.32432f
C302 3_OTA_0.OTA_stage1_0.vd2.t5 VGND 1.32432f
C303 3_OTA_0.OTA_stage1_0.vd2.t7 VGND 1.31571f
C304 3_OTA_0.OTA_stage1_0.vd2.t1 VGND 0.354781f
C305 3_OTA_0.OTA_stage1_0.vd2.t3 VGND 0.033828f
C306 3_OTA_0.OTA_stage1_0.vd2.t2 VGND 0.033816f
C307 3_OTA_0.3rd_3_OTA_0.vd4.n0 VGND 0.593328f
C308 3_OTA_0.3rd_3_OTA_0.vd4.n1 VGND 1.19513f
C309 3_OTA_0.3rd_3_OTA_0.vd4.t10 VGND 0.557947f
C310 3_OTA_0.3rd_3_OTA_0.vd4.t12 VGND 0.559799f
C311 3_OTA_0.3rd_3_OTA_0.vd4.n2 VGND 0.604581f
C312 3_OTA_0.3rd_3_OTA_0.vd4.t11 VGND 0.559799f
C313 3_OTA_0.3rd_3_OTA_0.vd4.t8 VGND 0.555128f
C314 3_OTA_0.3rd_3_OTA_0.vd4.t9 VGND 16.543098f
C315 3_OTA_0.3rd_3_OTA_0.vd4.t4 VGND 0.04967f
C316 3_OTA_0.3rd_3_OTA_0.vd4.t0 VGND 0.091357f
C317 3_OTA_0.3rd_3_OTA_0.vd4.t1 VGND 0.091357f
C318 3_OTA_0.3rd_3_OTA_0.vd4.n3 VGND 0.253746f
C319 3_OTA_0.3rd_3_OTA_0.vd4.t2 VGND 0.43452f
C320 3_OTA_0.3rd_3_OTA_0.vd4.t3 VGND 0.482932f
C321 3_OTA_0.3rd_3_OTA_0.vd4.n4 VGND 2.53677f
C322 3_OTA_0.3rd_3_OTA_0.vd4.n5 VGND 1.47312f
C323 3_OTA_0.3rd_3_OTA_0.vd4.n6 VGND 1.4592f
C324 3_OTA_0.3rd_3_OTA_0.vd4.t5 VGND 0.044809f
C325 3_OTA_0.3rd_3_OTA_0.vd4.t7 VGND 0.009136f
C326 3_OTA_0.3rd_3_OTA_0.vd4.t6 VGND 0.009136f
C327 3_OTA_0.3rd_3_OTA_0.vd4.n7 VGND 0.054041f
C328 a_12564_25551.t9 VGND 0.101734f
C329 a_12564_25551.t11 VGND 0.429436f
C330 a_12564_25551.t8 VGND 0.401468f
C331 a_12564_25551.t2 VGND 0.218001f
C332 a_12564_25551.t1 VGND 0.218001f
C333 a_12564_25551.n0 VGND 0.674641f
C334 a_12564_25551.t6 VGND 0.218001f
C335 a_12564_25551.t5 VGND 0.218001f
C336 a_12564_25551.n1 VGND 0.765785f
C337 a_12564_25551.n2 VGND 4.74835f
C338 a_12564_25551.t0 VGND 0.218001f
C339 a_12564_25551.t4 VGND 0.218001f
C340 a_12564_25551.n3 VGND 0.67477f
C341 a_12564_25551.t3 VGND 0.218001f
C342 a_12564_25551.t7 VGND 0.218001f
C343 a_12564_25551.n4 VGND 0.765807f
C344 a_12564_25551.n5 VGND 3.55783f
C345 a_12564_25551.n6 VGND 2.90218f
C346 a_12564_25551.n7 VGND 1.41326f
C347 a_12564_25551.n8 VGND 2.08198f
C348 a_12564_25551.n9 VGND 0.237014f
C349 a_12564_25551.t10 VGND 0.101734f
C350 3_OTA_0.OTA_vref_0.vb1.n0 VGND 5.75346f
C351 3_OTA_0.OTA_vref_0.vb1.n1 VGND 0.352136f
C352 3_OTA_0.OTA_vref_0.vb1.t9 VGND 0.858318f
C353 3_OTA_0.OTA_vref_0.vb1.t7 VGND 0.846486f
C354 3_OTA_0.OTA_vref_0.vb1.t8 VGND 0.846486f
C355 3_OTA_0.OTA_vref_0.vb1.t6 VGND 0.846486f
C356 3_OTA_0.OTA_vref_0.vb1.t0 VGND 0.007035f
C357 3_OTA_0.OTA_vref_0.vb1.t3 VGND 0.007035f
C358 3_OTA_0.OTA_vref_0.vb1.n2 VGND 0.018857f
C359 3_OTA_0.OTA_vref_0.vb1.t5 VGND 0.007035f
C360 3_OTA_0.OTA_vref_0.vb1.t4 VGND 0.007035f
C361 3_OTA_0.OTA_vref_0.vb1.n3 VGND 0.017824f
C362 3_OTA_0.OTA_vref_0.vb1.t2 VGND 0.007035f
C363 3_OTA_0.OTA_vref_0.vb1.t1 VGND 0.007035f
C364 3_OTA_0.OTA_vref_0.vb1.n4 VGND 0.017824f
C365 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n0 VGND 1.10559f
C366 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t0 VGND 0.076807f
C367 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t4 VGND 0.079082f
C368 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t26 VGND 0.079082f
C369 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n1 VGND 0.26329f
C370 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t14 VGND 0.079082f
C371 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t8 VGND 0.079082f
C372 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n2 VGND 0.253461f
C373 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n3 VGND 1.60391f
C374 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t3 VGND 0.079082f
C375 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t27 VGND 0.079082f
C376 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n4 VGND 0.253461f
C377 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n5 VGND 0.930699f
C378 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t24 VGND 0.079082f
C379 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t1 VGND 0.079082f
C380 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n6 VGND 0.253461f
C381 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n7 VGND 0.930699f
C382 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t6 VGND 0.079082f
C383 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t28 VGND 0.079082f
C384 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n8 VGND 0.253461f
C385 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n9 VGND 0.930699f
C386 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t23 VGND 0.079082f
C387 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t9 VGND 0.079082f
C388 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n10 VGND 0.253461f
C389 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n11 VGND 0.907084f
C390 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t17 VGND 0.079082f
C391 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t13 VGND 0.079082f
C392 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n12 VGND 0.277022f
C393 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t30 VGND 0.079082f
C394 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t21 VGND 0.079082f
C395 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n13 VGND 0.253461f
C396 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n14 VGND 1.70869f
C397 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t18 VGND 0.079082f
C398 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t5 VGND 0.079082f
C399 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n15 VGND 0.253461f
C400 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n16 VGND 0.921182f
C401 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t2 VGND 0.079082f
C402 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t16 VGND 0.079082f
C403 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n17 VGND 0.253461f
C404 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n18 VGND 0.921182f
C405 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t19 VGND 0.079082f
C406 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t10 VGND 0.079082f
C407 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n19 VGND 0.253461f
C408 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n20 VGND 0.921182f
C409 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t31 VGND 0.079082f
C410 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t15 VGND 0.079082f
C411 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n21 VGND 0.253461f
C412 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n22 VGND 0.921182f
C413 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t20 VGND 0.079082f
C414 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t12 VGND 0.079082f
C415 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n23 VGND 0.253461f
C416 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n24 VGND 0.921182f
C417 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t32 VGND 0.079082f
C418 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t25 VGND 0.079082f
C419 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n25 VGND 0.253461f
C420 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n26 VGND 1.42732f
C421 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t22 VGND 0.079082f
C422 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t11 VGND 0.079082f
C423 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n27 VGND 0.253331f
C424 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n28 VGND 1.30826f
C425 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t7 VGND 0.079082f
C426 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.t29 VGND 0.079082f
C427 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0.n29 VGND 0.253461f
C428 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 VGND 0.072231f
C429 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 VGND 0.110183f
C430 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 VGND 0.109159f
C431 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 VGND -3.71022f
C432 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 VGND 3.98508f
C433 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 VGND 0.480217f
C434 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 VGND 0.478981f
C435 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 VGND 1.17118f
C436 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 VGND 0.305431f
C437 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 VGND 0.478028f
C438 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 VGND 0.234187f
C439 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 VGND 0.470573f
C440 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 VGND 0.478028f
C441 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 VGND 0.470573f
C442 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 VGND 0.478028f
C443 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 VGND 0.470129f
C444 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 VGND 0.478028f
C445 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 VGND 0.119324f
C446 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 VGND 0.391163f
C447 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 VGND 0.207754f
C448 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 VGND 0.305316f
C449 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 VGND 0.478809f
C450 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 VGND 0.222027f
C451 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 VGND 0.474153f
C452 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 VGND 0.478028f
C453 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 VGND 0.474153f
C454 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 VGND 0.478028f
C455 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 VGND 0.472108f
C456 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 VGND 0.478028f
C457 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 VGND 0.114607f
C458 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 VGND 0.358209f
C459 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 VGND 0.171144f
C460 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 VGND 0.305164f
C461 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 VGND 0.478028f
C462 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 VGND 0.234725f
C463 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 VGND 0.471116f
C464 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 VGND 0.478028f
C465 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 VGND 0.471116f
C466 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 VGND 0.478028f
C467 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 VGND 0.471016f
C468 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 VGND 0.478028f
C469 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 VGND 0.116651f
C470 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 VGND 0.391917f
C471 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 VGND 0.175402f
C472 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 VGND 0.305187f
C473 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 VGND 0.478881f
C474 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 VGND 0.232796f
C475 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 VGND 0.470031f
C476 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 VGND 0.478028f
C477 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 VGND 0.470031f
C478 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 VGND 0.478028f
C479 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 VGND 0.470335f
C480 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 VGND 0.478028f
C481 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 VGND 0.118954f
C482 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 VGND 0.357235f
C483 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 VGND 0.171379f
C484 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 VGND 0.305728f
C485 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 VGND 0.478028f
C486 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 VGND 0.231521f
C487 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 VGND 0.470852f
C488 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 VGND 0.478028f
C489 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 VGND 0.470852f
C490 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 VGND 0.478028f
C491 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 VGND 0.466741f
C492 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 VGND 0.478028f
C493 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 VGND 0.124091f
C494 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 VGND 0.391922f
C495 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 VGND 0.175402f
C496 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 VGND 0.478028f
C497 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 VGND 0.282649f
C498 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 VGND 0.46793f
C499 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 VGND 0.478028f
C500 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 VGND 0.240285f
C501 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 VGND 0.478028f
C502 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 VGND 0.46793f
C503 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 VGND 0.304748f
C504 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 VGND 0.478028f
C505 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 VGND 0.303892f
C506 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 VGND 0.157746f
C507 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 VGND 0.205145f
C508 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 VGND 0.171854f
C509 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 VGND 0.305508f
C510 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 VGND 0.478028f
C511 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 VGND 0.22844f
C512 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 VGND 0.473853f
C513 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 VGND 0.478028f
C514 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 VGND 0.473853f
C515 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 VGND 0.478028f
C516 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 VGND 0.473079f
C517 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 VGND 0.478028f
C518 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 VGND 0.113695f
C519 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 VGND 0.395354f
C520 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 VGND 0.17643f
C521 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 VGND 0.480413f
C522 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 VGND 0.478986f
C523 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 VGND 1.18519f
C524 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 VGND 0.383039f
C525 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 VGND 0.473185f
C526 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 VGND 0.147422f
C527 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 VGND 0.215214f
C528 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 VGND 0.041255f
C529 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 VGND 0.04125f
C530 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 VGND 1.0568f
C531 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 VGND 0.444711f
C532 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 VGND 0.201225f
C533 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 VGND 0.215214f
C534 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 VGND 0.184059f
C535 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 VGND 0.10796f
C536 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 VGND 0.122425f
C537 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 VGND 0.110183f
C538 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 VGND 0.122425f
C539 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 VGND 0.490623f
C540 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 VGND 0.201231f
C541 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 VGND 0.381488f
C542 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 VGND 0.215214f
C543 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 VGND 0.329195f
C544 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 VGND 0.122425f
C545 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 VGND 0.21592f
C546 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 VGND 0.21592f
C547 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 VGND 0.101613f
C548 a_3013_4521.n0 VGND 0.297561f
C549 a_3013_4521.n1 VGND 0.29688f
C550 a_3013_4521.n2 VGND 0.297638f
C551 a_3013_4521.n3 VGND 0.2952f
C552 a_3013_4521.n4 VGND 0.5851f
C553 a_3013_4521.n5 VGND 0.294579f
C554 a_3013_4521.n6 VGND 0.296855f
C555 a_3013_4521.n7 VGND 0.755178f
C556 a_3013_4521.n8 VGND 0.296085f
C557 a_3013_4521.n9 VGND 0.293416f
C558 a_3013_4521.n10 VGND 0.294606f
C559 a_3013_4521.n11 VGND 0.292443f
C560 a_3013_4521.n12 VGND 0.23217f
C561 a_3013_4521.t9 VGND 0.036645f
C562 a_3013_4521.t28 VGND 0.036645f
C563 a_3013_4521.t0 VGND 0.036645f
C564 a_3013_4521.n13 VGND 0.078229f
C565 a_3013_4521.n14 VGND 0.188481f
C566 a_3013_4521.t43 VGND 0.428029f
C567 a_3013_4521.n15 VGND 0.126525f
C568 a_3013_4521.n16 VGND 0.13857f
C569 a_3013_4521.t35 VGND 0.428675f
C570 a_3013_4521.n17 VGND 0.188077f
C571 a_3013_4521.n18 VGND 0.174451f
C572 a_3013_4521.n19 VGND 0.188077f
C573 a_3013_4521.t27 VGND 0.428029f
C574 a_3013_4521.n20 VGND 0.191672f
C575 a_3013_4521.t7 VGND 0.036645f
C576 a_3013_4521.t34 VGND 0.036645f
C577 a_3013_4521.n21 VGND 0.078439f
C578 a_3013_4521.n22 VGND 0.109754f
C579 a_3013_4521.t17 VGND 0.428668f
C580 a_3013_4521.n23 VGND 0.499869f
C581 a_3013_4521.n24 VGND 0.184946f
C582 a_3013_4521.n25 VGND 0.126511f
C583 a_3013_4521.t29 VGND 0.428029f
C584 a_3013_4521.t18 VGND 0.036645f
C585 a_3013_4521.t47 VGND 0.036645f
C586 a_3013_4521.n26 VGND 0.078282f
C587 a_3013_4521.n27 VGND 0.280854f
C588 a_3013_4521.t10 VGND 0.036645f
C589 a_3013_4521.t30 VGND 0.036645f
C590 a_3013_4521.n28 VGND 0.078282f
C591 a_3013_4521.t12 VGND 0.036645f
C592 a_3013_4521.t22 VGND 0.036645f
C593 a_3013_4521.n29 VGND 0.078282f
C594 a_3013_4521.t40 VGND 0.036645f
C595 a_3013_4521.t2 VGND 0.036645f
C596 a_3013_4521.n30 VGND 0.078282f
C597 a_3013_4521.n31 VGND 0.224396f
C598 a_3013_4521.n32 VGND 0.074163f
C599 a_3013_4521.n33 VGND 0.12649f
C600 a_3013_4521.n34 VGND 0.19551f
C601 a_3013_4521.n35 VGND 0.194486f
C602 a_3013_4521.t39 VGND 0.428029f
C603 a_3013_4521.n36 VGND 0.234826f
C604 a_3013_4521.n37 VGND 0.160406f
C605 a_3013_4521.n38 VGND 0.27505f
C606 a_3013_4521.n39 VGND 0.252051f
C607 a_3013_4521.n40 VGND 0.127924f
C608 a_3013_4521.n41 VGND 0.190285f
C609 a_3013_4521.t33 VGND 0.428029f
C610 a_3013_4521.n42 VGND 0.194221f
C611 a_3013_4521.t19 VGND 0.428029f
C612 a_3013_4521.n43 VGND 0.192537f
C613 a_3013_4521.n44 VGND 0.126525f
C614 a_3013_4521.t20 VGND 0.036645f
C615 a_3013_4521.t4 VGND 0.036645f
C616 a_3013_4521.n45 VGND 0.078229f
C617 a_3013_4521.t1 VGND 0.036645f
C618 a_3013_4521.t38 VGND 0.036645f
C619 a_3013_4521.n46 VGND 0.078229f
C620 a_3013_4521.n47 VGND 0.251476f
C621 a_3013_4521.n48 VGND 0.133677f
C622 a_3013_4521.n49 VGND 0.192784f
C623 a_3013_4521.t37 VGND 0.428029f
C624 a_3013_4521.n50 VGND 0.196603f
C625 a_3013_4521.t31 VGND 0.428029f
C626 a_3013_4521.n51 VGND 0.19224f
C627 a_3013_4521.n52 VGND 0.126525f
C628 a_3013_4521.t32 VGND 0.036645f
C629 a_3013_4521.t45 VGND 0.036645f
C630 a_3013_4521.n53 VGND 0.078229f
C631 a_3013_4521.t3 VGND 0.036645f
C632 a_3013_4521.t42 VGND 0.036645f
C633 a_3013_4521.n54 VGND 0.078229f
C634 a_3013_4521.t41 VGND 0.428029f
C635 a_3013_4521.n55 VGND 0.192525f
C636 a_3013_4521.n56 VGND 0.12649f
C637 a_3013_4521.n57 VGND 0.126526f
C638 a_3013_4521.n58 VGND 0.252068f
C639 a_3013_4521.n59 VGND 0.174451f
C640 a_3013_4521.n60 VGND 0.160431f
C641 a_3013_4521.n61 VGND 0.116428f
C642 a_3013_4521.n62 VGND 0.191094f
C643 a_3013_4521.t21 VGND 0.428029f
C644 a_3013_4521.n63 VGND 0.181626f
C645 a_3013_4521.t15 VGND 0.428029f
C646 a_3013_4521.n64 VGND 0.11634f
C647 a_3013_4521.n65 VGND 0.0753f
C648 a_3013_4521.t16 VGND 0.036645f
C649 a_3013_4521.t5 VGND 0.036645f
C650 a_3013_4521.n66 VGND 0.078283f
C651 a_3013_4521.n67 VGND 0.22423f
C652 a_3013_4521.t11 VGND 0.036645f
C653 a_3013_4521.t24 VGND 0.036645f
C654 a_3013_4521.n68 VGND 0.078282f
C655 a_3013_4521.n69 VGND 0.210449f
C656 a_3013_4521.n70 VGND 0.152363f
C657 a_3013_4521.n71 VGND 0.209679f
C658 a_3013_4521.t23 VGND 0.428029f
C659 a_3013_4521.n72 VGND 0.197958f
C660 a_3013_4521.t13 VGND 0.428029f
C661 a_3013_4521.n73 VGND 0.222906f
C662 a_3013_4521.n74 VGND 0.152378f
C663 a_3013_4521.t14 VGND 0.036645f
C664 a_3013_4521.t46 VGND 0.036645f
C665 a_3013_4521.n75 VGND 0.078282f
C666 a_3013_4521.t6 VGND 0.036645f
C667 a_3013_4521.t36 VGND 0.036645f
C668 a_3013_4521.n76 VGND 0.078282f
C669 a_3013_4521.t26 VGND 0.036645f
C670 a_3013_4521.t8 VGND 0.036645f
C671 a_3013_4521.n77 VGND 0.078229f
C672 a_3013_4521.n78 VGND 0.501476f
C673 a_3013_4521.n79 VGND 0.213011f
C674 a_3013_4521.n80 VGND 0.230335f
C675 a_3013_4521.t25 VGND 0.428029f
C676 a_3013_4521.n81 VGND 0.191545f
C677 a_3013_4521.n82 VGND 0.191539f
C678 a_3013_4521.n83 VGND 0.12649f
C679 a_3013_4521.n84 VGND 0.078229f
C680 a_3013_4521.t44 VGND 0.036645f
C681 3_OTA_0.OTA_stage1_0.vd1.t1 VGND 1.59305f
C682 3_OTA_0.OTA_stage1_0.vd1.t3 VGND 1.6036f
C683 3_OTA_0.OTA_stage1_0.vd1.t2 VGND 1.6036f
C684 3_OTA_0.OTA_stage1_0.vd1.t0 VGND 1.59305f
C685 a_24889_22946.t1 VGND 26.271801f
C686 a_24889_22946.t0 VGND 0.028206f
C687 VDPWR.t56 VGND 0.007391f
C688 VDPWR.n0 VGND 0.086893f
C689 VDPWR.t62 VGND 0.007391f
C690 VDPWR.t60 VGND 0.001972f
C691 VDPWR.t54 VGND 0.001972f
C692 VDPWR.n1 VGND 0.004206f
C693 VDPWR.n2 VGND 0.259396f
C694 VDPWR.n3 VGND 0.074565f
C695 VDPWR.t49 VGND 9.86e-19
C696 VDPWR.t50 VGND 9.86e-19
C697 VDPWR.n4 VGND 0.002065f
C698 VDPWR.n5 VGND 0.080859f
C699 VDPWR.n6 VGND 0.146284f
C700 VDPWR.n7 VGND 0.096028f
C701 VDPWR.n8 VGND 0.14239f
C702 VDPWR.n9 VGND 0.096714f
C703 VDPWR.n10 VGND 0.038455f
C704 VDPWR.t48 VGND 0.110613f
C705 VDPWR.n11 VGND 0.153074f
C706 VDPWR.n12 VGND 0.022082f
C707 VDPWR.n13 VGND 0.060739f
C708 VDPWR.n14 VGND 0.014117f
C709 VDPWR.t61 VGND 0.156764f
C710 VDPWR.n15 VGND 0.023902f
C711 VDPWR.n16 VGND 0.095277f
C712 VDPWR.n17 VGND 0.107421f
C713 VDPWR.n18 VGND 0.107421f
C714 VDPWR.n19 VGND 0.025556f
C715 VDPWR.t63 VGND 0.007432f
C716 VDPWR.n20 VGND 0.280203f
C717 VDPWR.t58 VGND 0.007391f
C718 VDPWR.t52 VGND 0.007391f
C719 VDPWR.n21 VGND 0.120361f
C720 VDPWR.n22 VGND 0.134038f
C721 VDPWR.n23 VGND 0.278048f
C722 VDPWR.n24 VGND 0.15407f
C723 VDPWR.n25 VGND 0.062066f
C724 VDPWR.n26 VGND 0.107421f
C725 VDPWR.n27 VGND 0.107421f
C726 VDPWR.n28 VGND 0.103712f
C727 VDPWR.n29 VGND 0.086248f
C728 VDPWR.n30 VGND 0.020502f
C729 VDPWR.n31 VGND 0.020502f
C730 VDPWR.n32 VGND 0.246703f
C731 VDPWR.n33 VGND 0.188552f
C732 VDPWR.n35 VGND 0.135467f
C733 VDPWR.t51 VGND 0.129382f
C734 VDPWR.n36 VGND 0.179702f
C735 VDPWR.n37 VGND 0.042763f
C736 VDPWR.n38 VGND 0.184486f
C737 VDPWR.n39 VGND 0.176697f
C738 VDPWR.n40 VGND 0.115694f
C739 VDPWR.n41 VGND 0.041422f
C740 VDPWR.n42 VGND 0.014117f
C741 VDPWR.t57 VGND 0.156764f
C742 VDPWR.n45 VGND 0.014117f
C743 VDPWR.n46 VGND 0.174593f
C744 VDPWR.n47 VGND 0.174763f
C745 VDPWR.n48 VGND 0.061122f
C746 VDPWR.n49 VGND 0.014117f
C747 VDPWR.t55 VGND 0.156764f
C748 VDPWR.n52 VGND 0.014117f
C749 VDPWR.n53 VGND 0.061824f
C750 VDPWR.n54 VGND 0.172038f
C751 VDPWR.n55 VGND 0.17064f
C752 VDPWR.n56 VGND 0.025005f
C753 VDPWR.n58 VGND 0.107423f
C754 VDPWR.n59 VGND 0.014117f
C755 VDPWR.n61 VGND 0.107421f
C756 VDPWR.n62 VGND 0.096991f
C757 VDPWR.n63 VGND 0.115502f
C758 VDPWR.n64 VGND 0.064657f
C759 VDPWR.n65 VGND 0.011562f
C760 VDPWR.n66 VGND 0.230539f
C761 VDPWR.n67 VGND 0.027737f
C762 VDPWR.n68 VGND 0.03107f
C763 VDPWR.n69 VGND 0.023257f
C764 VDPWR.n70 VGND 0.023257f
C765 VDPWR.n71 VGND 0.035264f
C766 VDPWR.t59 VGND 0.079886f
C767 VDPWR.t53 VGND 0.114508f
C768 VDPWR.n72 VGND 0.126126f
C769 VDPWR.n73 VGND 0.060041f
C770 VDPWR.n74 VGND 0.188078f
C771 VDPWR.n75 VGND 0.066681f
C772 VDPWR.n76 VGND 0.135211f
C773 VDPWR.n77 VGND 0.049457f
C774 VDPWR.n78 VGND 0.051562f
C775 VDPWR.n79 VGND 0.076026f
C776 VDPWR.n80 VGND 0.1361f
C777 VDPWR.n81 VGND 0.039113f
C778 VDPWR.n82 VGND 1.51143f
C779 VDPWR.n83 VGND 2.60059f
C780 VDPWR.t23 VGND 0.003549f
C781 VDPWR.t20 VGND 0.003549f
C782 VDPWR.n84 VGND 0.007787f
C783 VDPWR.t24 VGND 0.003549f
C784 VDPWR.t21 VGND 0.003549f
C785 VDPWR.n85 VGND 0.007415f
C786 VDPWR.n86 VGND 0.08229f
C787 VDPWR.n87 VGND 0.55026f
C788 VDPWR.n88 VGND 0.394582f
C789 VDPWR.n89 VGND 0.10508f
C790 VDPWR.n90 VGND 0.10508f
C791 VDPWR.n91 VGND 0.724406f
C792 VDPWR.n92 VGND 1.24787f
C793 VDPWR.t22 VGND 1.95792f
C794 VDPWR.n93 VGND 1.83412f
C795 VDPWR.t19 VGND 1.95766f
C796 VDPWR.n94 VGND 1.24612f
C797 VDPWR.n95 VGND 0.780436f
C798 VDPWR.n96 VGND 0.697352f
C799 VDPWR.n97 VGND 0.936649f
C800 VDPWR.n98 VGND 0.553356f
C801 VDPWR.n99 VGND 1.0141f
C802 VDPWR.n100 VGND 0.233334f
C803 VDPWR.n101 VGND 0.364675f
C804 VDPWR.n102 VGND 0.241506f
C805 VDPWR.n103 VGND 0.645414f
C806 VDPWR.n104 VGND 0.115644f
C807 VDPWR.n105 VGND 0.115621f
C808 VDPWR.n106 VGND 0.527319f
C809 VDPWR.n107 VGND 0.004543f
C810 VDPWR.n108 VGND 0.067353f
C811 VDPWR.n109 VGND 0.065816f
C812 VDPWR.n110 VGND 0.210244f
C813 VDPWR.n111 VGND 0.164954f
C814 VDPWR.n112 VGND 0.24854f
C815 VDPWR.n113 VGND 0.41315f
C816 VDPWR.n114 VGND 0.125112f
C817 VDPWR.n115 VGND 0.416341f
C818 VDPWR.n116 VGND 0.00558f
C819 VDPWR.n117 VGND 0.095679f
C820 VDPWR.n118 VGND 0.744998f
C821 VDPWR.n119 VGND 0.297716f
C822 VDPWR.n120 VGND 0.297716f
C823 VDPWR.t44 VGND 0.475293f
C824 VDPWR.t68 VGND 0.391746f
C825 VDPWR.n121 VGND 0.324413f
C826 VDPWR.n122 VGND 0.223544f
C827 VDPWR.n123 VGND 0.184749f
C828 VDPWR.t45 VGND 0.013801f
C829 VDPWR.t69 VGND 0.013801f
C830 VDPWR.n124 VGND 0.03585f
C831 VDPWR.t14 VGND 0.013801f
C832 VDPWR.t26 VGND 0.013801f
C833 VDPWR.n125 VGND 0.035189f
C834 VDPWR.n126 VGND 0.563073f
C835 VDPWR.n127 VGND 0.111301f
C836 VDPWR.t67 VGND 0.004929f
C837 VDPWR.t46 VGND 0.004929f
C838 VDPWR.n128 VGND 0.010682f
C839 VDPWR.n129 VGND 0.333225f
C840 VDPWR.n130 VGND 0.317993f
C841 VDPWR.n131 VGND 0.839293f
C842 VDPWR.n132 VGND 1.27048f
C843 VDPWR.n133 VGND 0.008701f
C844 VDPWR.n134 VGND 0.102676f
C845 VDPWR.t28 VGND 0.004929f
C846 VDPWR.t47 VGND 0.004929f
C847 VDPWR.n135 VGND 0.010726f
C848 VDPWR.t12 VGND 0.01965f
C849 VDPWR.t5 VGND 0.019492f
C850 VDPWR.n136 VGND 0.103023f
C851 VDPWR.n137 VGND 0.019654f
C852 VDPWR.n138 VGND 0.014276f
C853 VDPWR.n139 VGND 0.009115f
C854 VDPWR.t4 VGND 0.124707f
C855 VDPWR.n140 VGND 0.008842f
C856 VDPWR.n141 VGND 0.060247f
C857 VDPWR.n142 VGND 0.821577f
C858 VDPWR.t27 VGND 1.55382f
C859 VDPWR.t0 VGND 1.30894f
C860 VDPWR.t29 VGND 1.54603f
C861 VDPWR.t17 VGND 1.31721f
C862 VDPWR.n143 VGND 0.694616f
C863 VDPWR.n144 VGND 0.338206f
C864 VDPWR.t41 VGND 0.004929f
C865 VDPWR.t1 VGND 0.004929f
C866 VDPWR.n145 VGND 0.010682f
C867 VDPWR.n146 VGND 0.082057f
C868 VDPWR.n147 VGND 0.038673f
C869 VDPWR.n148 VGND 0.073879f
C870 VDPWR.n149 VGND 0.067822f
C871 VDPWR.n150 VGND 0.24168f
C872 VDPWR.n151 VGND 0.343208f
C873 VDPWR.n152 VGND 0.150373f
C874 VDPWR.n153 VGND 0.136893f
C875 VDPWR.n154 VGND 0.519146f
C876 VDPWR.n155 VGND 0.311414f
C877 VDPWR.n156 VGND 0.027738f
C878 VDPWR.n157 VGND 0.679302f
C879 VDPWR.n158 VGND 0.081596f
C880 VDPWR.n159 VGND 0.875382f
C881 VDPWR.n160 VGND 0.081573f
C882 VDPWR.n161 VGND 0.114606f
C883 VDPWR.n162 VGND 0.216012f
C884 VDPWR.n163 VGND 0.034916f
C885 VDPWR.n164 VGND 0.097519f
C886 VDPWR.n166 VGND 0.008842f
C887 VDPWR.n167 VGND 0.009115f
C888 VDPWR.n168 VGND 0.011926f
C889 VDPWR.n169 VGND 0.008842f
C890 VDPWR.n170 VGND 0.009235f
C891 VDPWR.n171 VGND 0.009454f
C892 VDPWR.n172 VGND 0.115933f
C893 VDPWR.t11 VGND 0.124707f
C894 VDPWR.n173 VGND 0.009115f
C895 VDPWR.n174 VGND 0.122296f
C896 VDPWR.n175 VGND 0.069435f
C897 VDPWR.n176 VGND 0.043325f
C898 VDPWR.n177 VGND 0.009115f
C899 VDPWR.n179 VGND 0.097519f
C900 VDPWR.n180 VGND 0.044163f
C901 VDPWR.n181 VGND 0.018295f
C902 VDPWR.n182 VGND 0.162093f
C903 VDPWR.n183 VGND 0.033964f
C904 VDPWR.n184 VGND 0.150784f
C905 VDPWR.n185 VGND 0.048323f
C906 VDPWR.t18 VGND 0.004929f
C907 VDPWR.t30 VGND 0.004929f
C908 VDPWR.n186 VGND 0.010726f
C909 VDPWR.n187 VGND 0.173527f
C910 VDPWR.n188 VGND 0.03655f
C911 VDPWR.n189 VGND 0.124937f
C912 VDPWR.n190 VGND 0.178311f
C913 VDPWR.n191 VGND 0.48554f
C914 VDPWR.n192 VGND 0.062297f
C915 VDPWR.n193 VGND 0.04062f
C916 VDPWR.n194 VGND 0.034758f
C917 VDPWR.n195 VGND 0.215099f
C918 VDPWR.n196 VGND 0.426675f
C919 VDPWR.n197 VGND 1.14014f
C920 VDPWR.n198 VGND 0.603077f
C921 VDPWR.n199 VGND 0.235436f
C922 VDPWR.n200 VGND 0.167402f
C923 VDPWR.n201 VGND 0.179565f
C924 VDPWR.n202 VGND 0.013698f
C925 VDPWR.n203 VGND 0.202527f
C926 VDPWR.n204 VGND 0.041955f
C927 VDPWR.t25 VGND 0.475293f
C928 VDPWR.t13 VGND 0.391746f
C929 VDPWR.n205 VGND 0.261164f
C930 VDPWR.n206 VGND 0.041955f
C931 VDPWR.n207 VGND 0.487891f
C932 VDPWR.n208 VGND 0.274603f
C933 VDPWR.n209 VGND 0.010138f
C934 VDPWR.n210 VGND 0.379229f
C935 VDPWR.n211 VGND 0.248014f
C936 VDPWR.n212 VGND 0.380534f
C937 VDPWR.n213 VGND 0.173304f
C938 VDPWR.n214 VGND 0.523979f
C939 VDPWR.n215 VGND 2.28671f
C940 VDPWR.t38 VGND 2.70794f
C941 VDPWR.t43 VGND 1.61944f
C942 VDPWR.n216 VGND 1.15524f
C943 VDPWR.t10 VGND 1.84627f
C944 VDPWR.t37 VGND 2.47999f
C945 VDPWR.n217 VGND 1.91858f
C946 VDPWR.n218 VGND 0.326926f
C947 VDPWR.n219 VGND 0.394925f
C948 VDPWR.n220 VGND 0.130408f
C949 VDPWR.n221 VGND 0.368178f
C950 VDPWR.n222 VGND 0.409466f
C951 VDPWR.n223 VGND 0.375712f
C952 VDPWR.n224 VGND 1.11008f
C953 VDPWR.n225 VGND 1.72495f
C954 VDPWR.n226 VGND 0.188457p
C955 VDPWR.n227 VGND 4.37804f
C956 VDPWR.n228 VGND 4.2993f
C957 VDPWR.n229 VGND 3.9687f
C958 VDPWR.n230 VGND 25.632599f
C959 VDPWR.n231 VGND 1.18124f
C960 VDPWR.n232 VGND 3.68578f
C961 VDPWR.n233 VGND 28.897902f
C962 VDPWR.n234 VGND 4.174049f
C963 VDPWR.n235 VGND 20.8463f
C964 VDPWR.t16 VGND 9.86e-19
C965 VDPWR.t66 VGND 9.86e-19
C966 VDPWR.n236 VGND 0.002065f
C967 VDPWR.n237 VGND 0.080859f
C968 VDPWR.n238 VGND 0.230817f
C969 VDPWR.n239 VGND 0.051512f
C970 VDPWR.t42 VGND 0.001972f
C971 VDPWR.t40 VGND 0.001972f
C972 VDPWR.n240 VGND 0.004206f
C973 VDPWR.t9 VGND 0.007391f
C974 VDPWR.t3 VGND 0.007391f
C975 VDPWR.t7 VGND 0.007391f
C976 VDPWR.n241 VGND 0.133983f
C977 VDPWR.t70 VGND 0.007391f
C978 VDPWR.n242 VGND 0.120361f
C979 VDPWR.t65 VGND 0.007432f
C980 VDPWR.n243 VGND 0.280149f
C981 VDPWR.n244 VGND 0.016683f
C982 VDPWR.n245 VGND 0.051652f
C983 VDPWR.n246 VGND 0.014117f
C984 VDPWR.t6 VGND 0.156764f
C985 VDPWR.n247 VGND 0.219263f
C986 VDPWR.n248 VGND 0.045548f
C987 VDPWR.n250 VGND 0.188552f
C988 VDPWR.n251 VGND 0.081688f
C989 VDPWR.n252 VGND 0.020502f
C990 VDPWR.n253 VGND 0.135467f
C991 VDPWR.t64 VGND 0.129382f
C992 VDPWR.n254 VGND 0.179702f
C993 VDPWR.n255 VGND 0.020502f
C994 VDPWR.n256 VGND 0.045101f
C995 VDPWR.n257 VGND 0.190124f
C996 VDPWR.n258 VGND 0.129995f
C997 VDPWR.n259 VGND 0.025556f
C998 VDPWR.n261 VGND 0.107421f
C999 VDPWR.n262 VGND 0.023902f
C1000 VDPWR.n263 VGND 0.072608f
C1001 VDPWR.n264 VGND 0.107421f
C1002 VDPWR.n265 VGND 0.107421f
C1003 VDPWR.n266 VGND 0.025005f
C1004 VDPWR.n267 VGND 0.112905f
C1005 VDPWR.n268 VGND 0.107423f
C1006 VDPWR.n269 VGND 0.107421f
C1007 VDPWR.n270 VGND 0.036257f
C1008 VDPWR.n271 VGND 0.014117f
C1009 VDPWR.t8 VGND 0.156764f
C1010 VDPWR.n274 VGND 0.014117f
C1011 VDPWR.n275 VGND 0.048871f
C1012 VDPWR.n276 VGND 0.15071f
C1013 VDPWR.n277 VGND 0.151812f
C1014 VDPWR.n278 VGND 0.049651f
C1015 VDPWR.n279 VGND 0.014117f
C1016 VDPWR.t2 VGND 0.156764f
C1017 VDPWR.n282 VGND 0.014117f
C1018 VDPWR.n283 VGND 0.048955f
C1019 VDPWR.n284 VGND 0.154435f
C1020 VDPWR.n285 VGND 0.138251f
C1021 VDPWR.n286 VGND 0.014117f
C1022 VDPWR.n288 VGND 0.107421f
C1023 VDPWR.n289 VGND 0.071071f
C1024 VDPWR.n290 VGND 0.049886f
C1025 VDPWR.n291 VGND 0.154027f
C1026 VDPWR.n292 VGND 0.278144f
C1027 VDPWR.n293 VGND 0.120295f
C1028 VDPWR.n294 VGND 0.09646f
C1029 VDPWR.n295 VGND 0.136638f
C1030 VDPWR.n296 VGND 0.075896f
C1031 VDPWR.n297 VGND 0.259398f
C1032 VDPWR.n298 VGND 0.14239f
C1033 VDPWR.n299 VGND 0.066679f
C1034 VDPWR.n300 VGND 0.023258f
C1035 VDPWR.n301 VGND 0.188088f
C1036 VDPWR.n302 VGND 0.113604f
C1037 VDPWR.n303 VGND 0.060061f
C1038 VDPWR.n304 VGND 0.038473f
C1039 VDPWR.n305 VGND 0.027754f
C1040 VDPWR.n306 VGND 0.031087f
C1041 VDPWR.n307 VGND 0.153091f
C1042 VDPWR.t15 VGND 0.110613f
C1043 VDPWR.n308 VGND 0.246685f
C1044 VDPWR.t39 VGND 0.065871f
C1045 VDPWR.n309 VGND 0.021183f
C1046 VDPWR.n310 VGND 0.028349f
C1047 VDPWR.n311 VGND 0.011635f
C1048 VDPWR.n312 VGND 0.096592f
C1049 VDPWR.n313 VGND 0.135224f
C1050 VDPWR.n314 VGND 0.049408f
C1051 VDPWR.n315 VGND 0.096127f
C1052 VDPWR.n316 VGND 0.090608f
C1053 VDPWR.n317 VGND 6.37875f
C1054 VDPWR.t35 VGND 0.003549f
C1055 VDPWR.t33 VGND 0.003549f
C1056 VDPWR.n318 VGND 0.007787f
C1057 VDPWR.t36 VGND 0.003549f
C1058 VDPWR.t32 VGND 0.003549f
C1059 VDPWR.n319 VGND 0.007415f
C1060 VDPWR.n320 VGND 0.08229f
C1061 VDPWR.n321 VGND 0.55026f
C1062 VDPWR.n322 VGND 0.394582f
C1063 VDPWR.n323 VGND 0.10508f
C1064 VDPWR.n324 VGND 0.10508f
C1065 VDPWR.n325 VGND 0.724406f
C1066 VDPWR.n326 VGND 1.24787f
C1067 VDPWR.t34 VGND 1.95792f
C1068 VDPWR.n327 VGND 1.83412f
C1069 VDPWR.t31 VGND 1.95766f
C1070 VDPWR.n328 VGND 1.24612f
C1071 VDPWR.n329 VGND 0.780436f
C1072 VDPWR.n330 VGND 0.697352f
C1073 VDPWR.n331 VGND 0.936649f
C1074 VDPWR.n332 VGND 0.745189f
C1075 VDPWR.n333 VGND 1.30519f
C1076 VDPWR.n334 VGND 21.8217f
C1077 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n0 VGND 1.12223f
C1078 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t0 VGND 0.077096f
C1079 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t13 VGND 0.07938f
C1080 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t22 VGND 0.07938f
C1081 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n1 VGND 0.264281f
C1082 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t28 VGND 0.07938f
C1083 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t11 VGND 0.07938f
C1084 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n2 VGND 0.254416f
C1085 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n3 VGND 1.60994f
C1086 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t10 VGND 0.07938f
C1087 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t27 VGND 0.07938f
C1088 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n4 VGND 0.254416f
C1089 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n5 VGND 0.934202f
C1090 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t23 VGND 0.07938f
C1091 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t7 VGND 0.07938f
C1092 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n6 VGND 0.254416f
C1093 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n7 VGND 0.934202f
C1094 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t3 VGND 0.07938f
C1095 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t32 VGND 0.07938f
C1096 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n8 VGND 0.254416f
C1097 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n9 VGND 0.934202f
C1098 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t25 VGND 0.07938f
C1099 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t6 VGND 0.07938f
C1100 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n10 VGND 0.254416f
C1101 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n11 VGND 0.910498f
C1102 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t26 VGND 0.07938f
C1103 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t8 VGND 0.07938f
C1104 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n12 VGND 0.278065f
C1105 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t4 VGND 0.07938f
C1106 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t17 VGND 0.07938f
C1107 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n13 VGND 0.254416f
C1108 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n14 VGND 1.71512f
C1109 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t19 VGND 0.07938f
C1110 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t2 VGND 0.07938f
C1111 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n15 VGND 0.254416f
C1112 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n16 VGND 0.92465f
C1113 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t16 VGND 0.07938f
C1114 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t24 VGND 0.07938f
C1115 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n17 VGND 0.254416f
C1116 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n18 VGND 0.92465f
C1117 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t20 VGND 0.07938f
C1118 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t14 VGND 0.07938f
C1119 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n19 VGND 0.254416f
C1120 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n20 VGND 0.92465f
C1121 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t15 VGND 0.07938f
C1122 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t29 VGND 0.07938f
C1123 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n21 VGND 0.254416f
C1124 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n22 VGND 0.92465f
C1125 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t18 VGND 0.07938f
C1126 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t1 VGND 0.07938f
C1127 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n23 VGND 0.254416f
C1128 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n24 VGND 0.92465f
C1129 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t5 VGND 0.07938f
C1130 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t21 VGND 0.07938f
C1131 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n25 VGND 0.254416f
C1132 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n26 VGND 1.43269f
C1133 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t30 VGND 0.07938f
C1134 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t12 VGND 0.07938f
C1135 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n27 VGND 0.254284f
C1136 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n28 VGND 1.31318f
C1137 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t9 VGND 0.07938f
C1138 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.t31 VGND 0.07938f
C1139 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0.n29 VGND 0.254416f
C1140 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n0 VGND 3.66925f
C1141 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n1 VGND 6.26673f
C1142 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n2 VGND 0.951247f
C1143 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n3 VGND 3.35899f
C1144 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t20 VGND 0.60782f
C1145 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t26 VGND 0.584499f
C1146 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n4 VGND 1.65263f
C1147 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t23 VGND 0.584499f
C1148 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n5 VGND 0.976322f
C1149 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t24 VGND 0.584499f
C1150 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n6 VGND 0.97502f
C1151 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t21 VGND 0.584499f
C1152 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t22 VGND 0.303436f
C1153 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t25 VGND 0.303436f
C1154 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t1 VGND 0.025841f
C1155 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t0 VGND 0.458739f
C1156 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t2 VGND 0.458739f
C1157 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t3 VGND 0.02587f
C1158 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t18 VGND 0.054748f
C1159 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t6 VGND 0.054748f
C1160 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n7 VGND 0.20797f
C1161 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t5 VGND 0.054748f
C1162 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t13 VGND 0.054748f
C1163 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n8 VGND 0.20797f
C1164 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t9 VGND 0.054748f
C1165 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t7 VGND 0.054748f
C1166 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n9 VGND 0.20797f
C1167 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t11 VGND 0.054748f
C1168 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t14 VGND 0.054748f
C1169 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n10 VGND 0.236203f
C1170 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t10 VGND 0.276061f
C1171 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t19 VGND 0.054748f
C1172 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t17 VGND 0.054748f
C1173 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n11 VGND 0.20797f
C1174 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t8 VGND 0.054748f
C1175 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t12 VGND 0.054748f
C1176 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n12 VGND 0.20797f
C1177 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t15 VGND 0.301381f
C1178 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t16 VGND 0.054748f
C1179 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.t4 VGND 0.054748f
C1180 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr.n13 VGND 0.20797f
C1181 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 VGND 0.072231f
C1182 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 VGND 0.110183f
C1183 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 VGND 0.109159f
C1184 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 VGND -3.71022f
C1185 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 VGND 3.98507f
C1186 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 VGND 0.478981f
C1187 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 VGND 0.480213f
C1188 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 VGND 1.17119f
C1189 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 VGND 0.305431f
C1190 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 VGND 0.478028f
C1191 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 VGND 0.234187f
C1192 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 VGND 0.470573f
C1193 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 VGND 0.478028f
C1194 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 VGND 0.470573f
C1195 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 VGND 0.478028f
C1196 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 VGND 0.470129f
C1197 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 VGND 0.478028f
C1198 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 VGND 0.119324f
C1199 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 VGND 0.391163f
C1200 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 VGND 0.207747f
C1201 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 VGND 0.305316f
C1202 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 VGND 0.478809f
C1203 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 VGND 0.222027f
C1204 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 VGND 0.474153f
C1205 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 VGND 0.478028f
C1206 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 VGND 0.474153f
C1207 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 VGND 0.478028f
C1208 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 VGND 0.472108f
C1209 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 VGND 0.478028f
C1210 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 VGND 0.114607f
C1211 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 VGND 0.358056f
C1212 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 VGND 0.1713f
C1213 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 VGND 0.305164f
C1214 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 VGND 0.478028f
C1215 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 VGND 0.234725f
C1216 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 VGND 0.471116f
C1217 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 VGND 0.478028f
C1218 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 VGND 0.471116f
C1219 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 VGND 0.478028f
C1220 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 VGND 0.471016f
C1221 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 VGND 0.478028f
C1222 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 VGND 0.116651f
C1223 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 VGND 0.391917f
C1224 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 VGND 0.175402f
C1225 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 VGND 0.305187f
C1226 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 VGND 0.478881f
C1227 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 VGND 0.232796f
C1228 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 VGND 0.470031f
C1229 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 VGND 0.478028f
C1230 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 VGND 0.470031f
C1231 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 VGND 0.478028f
C1232 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 VGND 0.470335f
C1233 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 VGND 0.478028f
C1234 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 VGND 0.118954f
C1235 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 VGND 0.357235f
C1236 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 VGND 0.171379f
C1237 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 VGND 0.305728f
C1238 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 VGND 0.478028f
C1239 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 VGND 0.231521f
C1240 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 VGND 0.470851f
C1241 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 VGND 0.478028f
C1242 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 VGND 0.470852f
C1243 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 VGND 0.478028f
C1244 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 VGND 0.466741f
C1245 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 VGND 0.478028f
C1246 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 VGND 0.124091f
C1247 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 VGND 0.391922f
C1248 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 VGND 0.175402f
C1249 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 VGND 0.478028f
C1250 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 VGND 0.28265f
C1251 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 VGND 0.46793f
C1252 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 VGND 0.478028f
C1253 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 VGND 0.240285f
C1254 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 VGND 0.478028f
C1255 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 VGND 0.46793f
C1256 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 VGND 0.304748f
C1257 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 VGND 0.478028f
C1258 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 VGND 0.303889f
C1259 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 VGND 0.157732f
C1260 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 VGND 0.205161f
C1261 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 VGND 0.171854f
C1262 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 VGND 0.305508f
C1263 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 VGND 0.478028f
C1264 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 VGND 0.22844f
C1265 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 VGND 0.473853f
C1266 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 VGND 0.478028f
C1267 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 VGND 0.473853f
C1268 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 VGND 0.478028f
C1269 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 VGND 0.473079f
C1270 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 VGND 0.478028f
C1271 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 VGND 0.113695f
C1272 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 VGND 0.395354f
C1273 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 VGND 0.17643f
C1274 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 VGND 0.480413f
C1275 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 VGND 0.478986f
C1276 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 VGND 1.18519f
C1277 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 VGND 0.383039f
C1278 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 VGND 0.473185f
C1279 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 VGND 0.215214f
C1280 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 VGND 0.201225f
C1281 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 VGND 0.215214f
C1282 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 VGND 0.215214f
C1283 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 VGND 0.184059f
C1284 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 VGND 0.04125f
C1285 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 VGND 0.041255f
C1286 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 VGND 1.0568f
C1287 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 VGND 0.444711f
C1288 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 VGND 0.122425f
C1289 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 VGND 0.110183f
C1290 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 VGND 0.10796f
C1291 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 VGND 0.122425f
C1292 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 VGND 0.490623f
C1293 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 VGND 0.201231f
C1294 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 VGND 0.381488f
C1295 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 VGND 0.147422f
C1296 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 VGND 0.329195f
C1297 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 VGND 0.122425f
C1298 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 VGND 0.21592f
C1299 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 VGND 0.21592f
C1300 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 VGND 0.101613f
C1301 a_12378_15906.n0 VGND 0.297823f
C1302 a_12378_15906.n1 VGND 0.297439f
C1303 a_12378_15906.n2 VGND 0.29823f
C1304 a_12378_15906.n3 VGND 0.29615f
C1305 a_12378_15906.n4 VGND 0.755844f
C1306 a_12378_15906.n5 VGND 0.585351f
C1307 a_12378_15906.n6 VGND 0.126637f
C1308 a_12378_15906.n7 VGND 0.297117f
C1309 a_12378_15906.n8 VGND 0.294839f
C1310 a_12378_15906.n9 VGND 0.295296f
C1311 a_12378_15906.n10 VGND 0.293675f
C1312 a_12378_15906.n11 VGND 0.295194f
C1313 a_12378_15906.n12 VGND 0.292701f
C1314 a_12378_15906.n13 VGND 0.160573f
C1315 a_12378_15906.n14 VGND 0.232375f
C1316 a_12378_15906.t41 VGND 0.036678f
C1317 a_12378_15906.n15 VGND 0.210635f
C1318 a_12378_15906.n16 VGND 0.152497f
C1319 a_12378_15906.n17 VGND 0.209864f
C1320 a_12378_15906.t22 VGND 0.428407f
C1321 a_12378_15906.n18 VGND 0.198133f
C1322 a_12378_15906.t16 VGND 0.428407f
C1323 a_12378_15906.t38 VGND 0.429053f
C1324 a_12378_15906.n19 VGND 0.501918f
C1325 a_12378_15906.n20 VGND 0.235053f
C1326 a_12378_15906.n21 VGND 0.188243f
C1327 a_12378_15906.t18 VGND 0.428407f
C1328 a_12378_15906.n22 VGND 0.191841f
C1329 a_12378_15906.t6 VGND 0.036678f
C1330 a_12378_15906.t11 VGND 0.036678f
C1331 a_12378_15906.n23 VGND 0.078298f
C1332 a_12378_15906.n24 VGND 0.188647f
C1333 a_12378_15906.t24 VGND 0.428407f
C1334 a_12378_15906.n25 VGND 0.126636f
C1335 a_12378_15906.n26 VGND 0.252394f
C1336 a_12378_15906.t10 VGND 0.428407f
C1337 a_12378_15906.n27 VGND 0.191714f
C1338 a_12378_15906.n28 VGND 0.191708f
C1339 a_12378_15906.n29 VGND 0.126601f
C1340 a_12378_15906.t25 VGND 0.036678f
C1341 a_12378_15906.t40 VGND 0.036678f
C1342 a_12378_15906.n30 VGND 0.078298f
C1343 a_12378_15906.t2 VGND 0.036678f
C1344 a_12378_15906.t19 VGND 0.036678f
C1345 a_12378_15906.n31 VGND 0.078298f
C1346 a_12378_15906.n32 VGND 0.190453f
C1347 a_12378_15906.t15 VGND 0.036678f
C1348 a_12378_15906.t47 VGND 0.036678f
C1349 a_12378_15906.n33 VGND 0.078298f
C1350 a_12378_15906.t4 VGND 0.036678f
C1351 a_12378_15906.t29 VGND 0.036678f
C1352 a_12378_15906.n34 VGND 0.078298f
C1353 a_12378_15906.t27 VGND 0.036678f
C1354 a_12378_15906.t46 VGND 0.036678f
C1355 a_12378_15906.n35 VGND 0.078508f
C1356 a_12378_15906.n36 VGND 0.109851f
C1357 a_12378_15906.n37 VGND 0.128037f
C1358 a_12378_15906.t26 VGND 0.428407f
C1359 a_12378_15906.n38 VGND 0.194392f
C1360 a_12378_15906.n39 VGND 0.192707f
C1361 a_12378_15906.t28 VGND 0.428407f
C1362 a_12378_15906.n40 VGND 0.252273f
C1363 a_12378_15906.n41 VGND 0.285147f
C1364 a_12378_15906.n42 VGND 0.185109f
C1365 a_12378_15906.n43 VGND 0.126622f
C1366 a_12378_15906.t20 VGND 0.428407f
C1367 a_12378_15906.t23 VGND 0.036678f
C1368 a_12378_15906.t3 VGND 0.036678f
C1369 a_12378_15906.n44 VGND 0.078351f
C1370 a_12378_15906.t1 VGND 0.036678f
C1371 a_12378_15906.t37 VGND 0.036678f
C1372 a_12378_15906.n45 VGND 0.078353f
C1373 a_12378_15906.n46 VGND 0.224428f
C1374 a_12378_15906.n47 VGND 0.075366f
C1375 a_12378_15906.n48 VGND 0.191262f
C1376 a_12378_15906.t32 VGND 0.428407f
C1377 a_12378_15906.n49 VGND 0.116443f
C1378 a_12378_15906.n50 VGND 0.188243f
C1379 a_12378_15906.t36 VGND 0.428407f
C1380 a_12378_15906.n51 VGND 0.181786f
C1381 a_12378_15906.n52 VGND 0.116531f
C1382 a_12378_15906.t33 VGND 0.036678f
C1383 a_12378_15906.t42 VGND 0.036678f
C1384 a_12378_15906.n53 VGND 0.078351f
C1385 a_12378_15906.t44 VGND 0.036678f
C1386 a_12378_15906.t9 VGND 0.036678f
C1387 a_12378_15906.n54 VGND 0.078351f
C1388 a_12378_15906.n55 VGND 0.224594f
C1389 a_12378_15906.n56 VGND 0.074228f
C1390 a_12378_15906.t34 VGND 0.429046f
C1391 a_12378_15906.n57 VGND 0.512311f
C1392 a_12378_15906.t5 VGND 0.036678f
C1393 a_12378_15906.t35 VGND 0.036678f
C1394 a_12378_15906.n58 VGND 0.078351f
C1395 a_12378_15906.n59 VGND 0.281102f
C1396 a_12378_15906.t21 VGND 0.036678f
C1397 a_12378_15906.t45 VGND 0.036678f
C1398 a_12378_15906.n60 VGND 0.078351f
C1399 a_12378_15906.n61 VGND 0.126601f
C1400 a_12378_15906.n62 VGND 0.195683f
C1401 a_12378_15906.n63 VGND 0.194658f
C1402 a_12378_15906.t8 VGND 0.428407f
C1403 a_12378_15906.n64 VGND 0.213178f
C1404 a_12378_15906.n65 VGND 0.138692f
C1405 a_12378_15906.n66 VGND 0.15275f
C1406 a_12378_15906.n67 VGND 0.229843f
C1407 a_12378_15906.n68 VGND 0.133795f
C1408 a_12378_15906.n69 VGND 0.192954f
C1409 a_12378_15906.t14 VGND 0.428407f
C1410 a_12378_15906.n70 VGND 0.196777f
C1411 a_12378_15906.t30 VGND 0.428407f
C1412 a_12378_15906.n71 VGND 0.19241f
C1413 a_12378_15906.n72 VGND 0.126637f
C1414 a_12378_15906.t0 VGND 0.036678f
C1415 a_12378_15906.t31 VGND 0.036678f
C1416 a_12378_15906.n73 VGND 0.078298f
C1417 a_12378_15906.t13 VGND 0.036678f
C1418 a_12378_15906.t43 VGND 0.036678f
C1419 a_12378_15906.n74 VGND 0.078298f
C1420 a_12378_15906.t12 VGND 0.428407f
C1421 a_12378_15906.n75 VGND 0.192695f
C1422 a_12378_15906.n76 VGND 0.126601f
C1423 a_12378_15906.n77 VGND 0.126638f
C1424 a_12378_15906.n78 VGND 0.230436f
C1425 a_12378_15906.n79 VGND 0.15275f
C1426 a_12378_15906.n80 VGND 0.160547f
C1427 a_12378_15906.n81 VGND 0.244957f
C1428 a_12378_15906.n82 VGND 0.152512f
C1429 a_12378_15906.t7 VGND 0.036678f
C1430 a_12378_15906.t17 VGND 0.036678f
C1431 a_12378_15906.n83 VGND 0.078351f
C1432 a_12378_15906.n84 VGND 0.078351f
C1433 a_12378_15906.t39 VGND 0.036678f
C1434 a_18163_10306.t0 VGND 23.3704f
C1435 a_18163_10306.n0 VGND 2.20167f
C1436 a_18163_10306.t1 VGND 0.029528f
C1437 a_18163_10306.t2 VGND 0.029518f
C1438 a_18163_10306.t3 VGND 0.233892f
C1439 a_18163_10306.t4 VGND 0.435024f
C1440 ua[2].t2 VGND 0.771754f
C1441 ua[2].t1 VGND 0.405603f
C1442 ua[2].n0 VGND 0.886904f
C1443 ua[2].t3 VGND 0.771752f
C1444 ua[2].t0 VGND 0.405603f
C1445 ua[2].n1 VGND 0.886906f
C1446 ua[2].n2 VGND 0.731678f
C1447 3_OTA_0.3rd_3_OTA_0.vd3.n0 VGND 0.456197f
C1448 3_OTA_0.3rd_3_OTA_0.vd3.n1 VGND 1.97994f
C1449 3_OTA_0.3rd_3_OTA_0.vd3.n2 VGND 1.83635f
C1450 3_OTA_0.3rd_3_OTA_0.vd3.n3 VGND 0.036861f
C1451 3_OTA_0.3rd_3_OTA_0.vd3.n4 VGND 1.84565f
C1452 3_OTA_0.3rd_3_OTA_0.vd3.n5 VGND 2.01844f
C1453 3_OTA_0.3rd_3_OTA_0.vd3.t14 VGND 0.292323f
C1454 3_OTA_0.3rd_3_OTA_0.vd3.t17 VGND 0.292237f
C1455 3_OTA_0.3rd_3_OTA_0.vd3.t16 VGND 0.292237f
C1456 3_OTA_0.3rd_3_OTA_0.vd3.t13 VGND 0.291885f
C1457 3_OTA_0.3rd_3_OTA_0.vd3.t1 VGND 0.047867f
C1458 3_OTA_0.3rd_3_OTA_0.vd3.t2 VGND 0.047867f
C1459 3_OTA_0.3rd_3_OTA_0.vd3.n6 VGND 0.150905f
C1460 3_OTA_0.3rd_3_OTA_0.vd3.t3 VGND 0.241422f
C1461 3_OTA_0.3rd_3_OTA_0.vd3.t0 VGND 0.218393f
C1462 3_OTA_0.3rd_3_OTA_0.vd3.n7 VGND 0.638972f
C1463 3_OTA_0.3rd_3_OTA_0.vd3.t5 VGND 0.016894f
C1464 3_OTA_0.3rd_3_OTA_0.vd3.t7 VGND 0.016894f
C1465 3_OTA_0.3rd_3_OTA_0.vd3.t6 VGND 0.665688f
C1466 3_OTA_0.3rd_3_OTA_0.vd3.t18 VGND 0.665686f
C1467 3_OTA_0.3rd_3_OTA_0.vd3.n8 VGND 0.248119f
C1468 3_OTA_0.3rd_3_OTA_0.vd3.t12 VGND 0.665688f
C1469 3_OTA_0.3rd_3_OTA_0.vd3.t10 VGND 0.665686f
C1470 3_OTA_0.3rd_3_OTA_0.vd3.n9 VGND 0.248119f
C1471 3_OTA_0.3rd_3_OTA_0.vd3.t11 VGND 0.004787f
C1472 3_OTA_0.3rd_3_OTA_0.vd3.t9 VGND 0.004787f
C1473 3_OTA_0.3rd_3_OTA_0.vd3.n10 VGND 0.010125f
C1474 3_OTA_0.3rd_3_OTA_0.vd3.t15 VGND 0.665688f
C1475 3_OTA_0.3rd_3_OTA_0.vd3.t8 VGND 0.665686f
C1476 3_OTA_0.3rd_3_OTA_0.vd3.n11 VGND 0.248119f
C1477 3_OTA_0.3rd_3_OTA_0.vd3.t4 VGND 0.665688f
C1478 3_OTA_0.3rd_3_OTA_0.vd3.t19 VGND 0.665686f
C1479 3_OTA_0.3rd_3_OTA_0.vd3.n12 VGND 0.248119f
C1480 3_OTA_0.3rd_3_OTA_0.vd3.n13 VGND 1.78256f
.ends

