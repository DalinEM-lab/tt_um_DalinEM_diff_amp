* NGSPICE file created from BGR_BJT_final_flat.ext - technology: sky130A

.subckt BGR_BJT_final_flat vcc vss vref
X0 BGR_BJT_stage1_0.vref0.t21 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 BGR_BJT_stage1_0.vr.t9 vss.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X1 vss.t26 a_365_2822.t30 a_365_2822.t31 vss.t25 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X2 a_2451_1374# a_2251_1286# BGR_BJT_stage1_0.vref0.t0 vss.t48 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X3 a_3741_1374# a_3541_1286# a_3541_1286# vss.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X4 a_365_2822.t47 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 BGR_BJT_stage1_0.vref0.t27 vss.t53 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X5 vss.t43 vss.t42 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X6 vcc.t17 BGR_BJT_stage1_0.vr.t2 BGR_BJT_stage1_0.vr.t3 vcc.t16 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=5800,316 d=2900,158
X7 a_365_2822.t46 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 BGR_BJT_stage1_0.vref0.t29 vss.t55 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X8 a_365_2822.t29 a_365_2822.t28 vss.t34 vss.t33 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X9 BGR_BJT_stage1_0.vr.t14 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 BGR_BJT_stage1_0.vref0.t20 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X10 a_365_2822.t45 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 BGR_BJT_stage1_0.vref0.t28 vss.t54 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X11 vss.t28 a_365_2822.t26 a_365_2822.t27 vss.t27 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X12 a_2251_1286# BGR_BJT_stage1_0.vr.t20 vcc.t7 vcc.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X13 a_4831_1286# BGR_BJT_stage1_0.vr.t21 vcc.t15 vcc.t14 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X14 a_365_2822.t44 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 BGR_BJT_stage1_0.vref0.t1 vss.t51 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X15 BGR_BJT_stage1_0.vref0.t19 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 BGR_BJT_stage1_0.vr.t16 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X16 a_365_2822.t43 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 BGR_BJT_stage1_0.vref0.t22 vss.t49 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X17 vss.t18 a_365_2822.t24 a_365_2822.t25 vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X18 BGR_BJT_stage1_0.vref0.t18 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 BGR_BJT_stage1_0.vr.t8 vss.t35 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X19 a_365_2822.t42 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 BGR_BJT_stage1_0.vref0.t26 vss.t43 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X20 BGR_BJT_stage1_0.vref0.t2 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 a_365_2822.t41 vss.t50 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X21 a_5031_1374# a_4831_1286# a_4831_1286# vss.t60 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X22 a_4831_1286# a_4831_1286# a_5031_1374# vss.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X23 BGR_BJT_stage1_0.vr.t1 BGR_BJT_stage1_0.vr.t0 vcc.t3 vcc.t2 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=2900,158 d=5800,316
X24 a_365_2822.t23 a_365_2822.t22 vss.t1 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X25 a_2251_1286# a_2251_1286# a_2451_1374# vss.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X26 a_4831_1286# a_4831_1286# a_5031_1374# vss.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X27 vref.t4 a_6121_1286# a_6121_1286# vss.t41 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=11600,516
X28 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 BGR_BJT_stage1_0.vr.t22 vcc.t13 vcc.t12 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=11600,516
X29 a_3541_1286# BGR_BJT_stage1_0.vr.t23 vcc.t11 vcc.t10 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X30 a_6121_1286# BGR_BJT_stage1_0.vr.t24 vcc.t9 vcc.t8 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X31 BGR_BJT_stage1_0.vref0.t17 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 BGR_BJT_stage1_0.vr.t18 vss.t23 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X32 vss.t30 a_365_2822.t20 a_365_2822.t21 vss.t29 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X33 BGR_BJT_stage1_0.vr.t11 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 BGR_BJT_stage1_0.vref0.t16 vss.t21 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X34 a_365_2822.t19 a_365_2822.t18 vss.t20 vss.t19 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X35 BGR_BJT_stage1_0.vref0.t23 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 a_365_2822.t40 vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X36 BGR_BJT_stage1_0.vref0.t15 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 BGR_BJT_stage1_0.vr.t6 vss.t31 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X37 vss.t5 a_365_2822.t16 a_365_2822.t17 vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X38 BGR_BJT_stage1_0.vref0.t25 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 a_365_2822.t39 vss.t55 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X39 BGR_BJT_stage1_0.vr.t17 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 BGR_BJT_stage1_0.vref0.t14 vss.t27 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X40 a_3541_1286# a_3541_1286# a_3741_1374# vss.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X41 a_5031_1374# a_4831_1286# a_4831_1286# vss.t57 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X42 BGR_BJT_stage1_0.vref0.t13 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 BGR_BJT_stage1_0.vr.t13 vss.t33 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X43 vss.t7 a_365_2822.t14 a_365_2822.t15 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X44 BGR_BJT_stage1_0.vref0.t3 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 a_365_2822.t38 vss.t54 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X45 a_2451_1374# a_2251_1286# a_2251_1286# vss.t46 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X46 a_3741_1374# a_3541_1286# a_2451_1374# vss.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X47 vcc.t5 BGR_BJT_stage1_0.vr.t25 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X48 BGR_BJT_stage1_0.vref0.t32 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 a_365_2822.t37 vss.t43 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X49 a_365_2822.t13 a_365_2822.t12 vss.t36 vss.t35 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X50 vss.t3 a_365_2822.t10 a_365_2822.t11 vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X51 a_365_2822.t9 a_365_2822.t8 vss.t9 vss.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X52 BGR_BJT_stage1_0.vr.t19 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 BGR_BJT_stage1_0.vref0.t12 vss.t25 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X53 BGR_BJT_stage1_0.vref0.t4 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 a_365_2822.t36 vss.t53 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X54 a_365_2822.t7 a_365_2822.t6 vss.t24 vss.t23 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X55 BGR_BJT_stage1_0.vr.t5 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 BGR_BJT_stage1_0.vref0.t11 vss.t29 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X56 a_365_2822.t35 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 BGR_BJT_stage1_0.vref0.t30 vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X57 vss.t22 a_365_2822.t4 a_365_2822.t5 vss.t21 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X58 a_365_2822.t3 a_365_2822.t2 vss.t32 vss.t31 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X59 BGR_BJT_stage1_0.vref0.t10 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 BGR_BJT_stage1_0.vr.t4 vss.t19 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X60 a_2251_1286# a_2251_1286# a_2451_1374# vss.t45 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X61 a_3541_1286# a_3541_1286# a_3741_1374# vss.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X62 a_6121_1286# a_6121_1286# vref.t3 vss.t40 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X63 vref.t2 a_6121_1286# a_6121_1286# vss.t39 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X64 a_3741_1374# a_3541_1286# a_3541_1286# vss.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X65 vref.t5 a_6121_1286# a_5031_1374# vss.t38 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X66 BGR_BJT_stage1_0.vr.t10 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 BGR_BJT_stage1_0.vref0.t9 vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X67 BGR_BJT_stage1_0.vref0.t5 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 a_365_2822.t34 vss.t51 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X68 a_365_2822.t1 a_365_2822.t0 vss.t11 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X69 BGR_BJT_stage1_0.vr.t12 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 BGR_BJT_stage1_0.vref0.t8 vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X70 a_365_2822.t33 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 BGR_BJT_stage1_0.vref0.t31 vss.t50 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X71 BGR_BJT_stage1_0.vref0.t24 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 a_365_2822.t32 vss.t49 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X72 vref.t0 BGR_BJT_stage1_0.vr.t26 vcc.t1 vcc.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X73 BGR_BJT_stage1_0.vref0.t7 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 BGR_BJT_stage1_0.vr.t15 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X74 BGR_BJT_stage1_0.vr.t7 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 BGR_BJT_stage1_0.vref0.t6 vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X75 a_2451_1374# a_2251_1286# a_2251_1286# vss.t44 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X76 a_5031_1374# a_4831_1286# a_3741_1374# vss.t56 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X77 a_6121_1286# a_6121_1286# vref.t1 vss.t37 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
R0 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 235.982
R1 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 235.978
R2 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 190.305
R3 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 190.305
R4 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 190.305
R5 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 190.305
R6 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 190.305
R7 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 190.305
R8 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 190.305
R9 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 190.305
R10 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 190.305
R11 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 190.305
R12 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 95.3656
R13 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 95.1789
R14 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 95.1648
R15 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 95.1535
R16 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 94.8416
R17 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 94.841
R18 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 94.8396
R19 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 94.8314
R20 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 94.8314
R21 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 94.8314
R22 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 94.8314
R23 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 94.8314
R24 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 94.8314
R25 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 94.8314
R26 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 94.8314
R27 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 94.8314
R28 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 94.8314
R29 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 94.8314
R30 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 94.8314
R31 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 94.8314
R32 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 94.8314
R33 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 94.8314
R34 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 94.8314
R35 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 94.8314
R36 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 94.8314
R37 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 94.8314
R38 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 94.8314
R39 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 83.7933
R40 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 83.5719
R41 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 83.5719
R42 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 83.5719
R43 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 83.5719
R44 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 73.3165
R45 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 26.074
R46 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 26.074
R47 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 26.074
R48 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 25.7843
R49 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 25.7843
R50 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 10.2824
R51 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 9.5389
R52 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 7.22993
R53 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 7.22993
R54 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 7.22993
R55 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 6.83022
R56 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 6.81633
R57 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 6.81633
R58 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 6.81633
R59 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 6.75312
R60 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 2.29815
R61 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 2.20008
R62 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 1.86108
R63 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 1.86108
R64 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 1.86108
R65 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 1.86108
R66 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 1.86108
R67 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 1.86108
R68 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 1.86108
R69 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 1.5505
R70 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 1.5505
R71 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 1.5505
R72 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 1.5505
R73 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 1.5505
R74 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 1.43912
R75 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 1.327
R76 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 1.32184
R77 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 1.27838
R78 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 1.26044
R79 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 1.24668
R80 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 1.19225
R81 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 1.1424
R82 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 1.11251
R83 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 1.10979
R84 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 1.10442
R85 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 1.10164
R86 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 1.10164
R87 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 1.10164
R88 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 1.10164
R89 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 1.10145
R90 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 1.09892
R91 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 1.09349
R92 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 1.09349
R93 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 1.08805
R94 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 1.08262
R95 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 1.08262
R96 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 1.08262
R97 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 1.07024
R98 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.959578
R99 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.885803
R100 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 0.77514
R101 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 0.756696
R102 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 0.679848
R103 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 0.645119
R104 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 0.645119
R105 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.645119
R106 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 0.645119
R107 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 0.645119
R108 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 0.645119
R109 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 0.645119
R110 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.645119
R111 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 0.645119
R112 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 0.645119
R113 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 0.645119
R114 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 0.645119
R115 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 0.645119
R116 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 0.645119
R117 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 0.645119
R118 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.645119
R119 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 0.645119
R120 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 0.645119
R121 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 0.645119
R122 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 0.645119
R123 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 0.645119
R124 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 0.645119
R125 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.645119
R126 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 0.645119
R127 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 0.645119
R128 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 0.645119
R129 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 0.628893
R130 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 0.628893
R131 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.590702
R132 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 0.570883
R133 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.498483
R134 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 0.495065
R135 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 0.495065
R136 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.481478
R137 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 0.481478
R138 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 0.475521
R139 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 0.470609
R140 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 0.470609
R141 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 0.465174
R142 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 0.465174
R143 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 0.465174
R144 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 0.459844
R145 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.459739
R146 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 0.459739
R147 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 0.446152
R148 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 0.446152
R149 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 0.445943
R150 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 0.443435
R151 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 0.440717
R152 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 0.434551
R153 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 0.414484
R154 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 0.408265
R155 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 0.408265
R156 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.406264
R157 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 0.40372
R158 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 0.40372
R159 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 0.290206
R160 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.0222391
R161 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 0.0209918
R162 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 0.0209918
R163 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 0.0209918
R164 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 0.0209918
R165 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 0.0183279
R166 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 0.00925374
R167 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 0.00730856
R168 BGR_BJT_stage1_0.vr.n0 BGR_BJT_stage1_0.vr.t3 651.943
R169 BGR_BJT_stage1_0.vr.n0 BGR_BJT_stage1_0.vr.t1 651.678
R170 BGR_BJT_stage1_0.vr.n0 BGR_BJT_stage1_0.vr.t25 60.1752
R171 BGR_BJT_stage1_0.vr.n0 BGR_BJT_stage1_0.vr.t22 60.088
R172 BGR_BJT_stage1_0.vr.n2 BGR_BJT_stage1_0.vr.t19 28.5589
R173 BGR_BJT_stage1_0.vr.n1 BGR_BJT_stage1_0.vr.t8 27.6016
R174 BGR_BJT_stage1_0.vr.n3 BGR_BJT_stage1_0.vr.t26 26.8562
R175 BGR_BJT_stage1_0.vr.n3 BGR_BJT_stage1_0.vr.t24 26.0492
R176 BGR_BJT_stage1_0.vr.n4 BGR_BJT_stage1_0.vr.t21 26.0492
R177 BGR_BJT_stage1_0.vr.n5 BGR_BJT_stage1_0.vr.t23 26.0492
R178 BGR_BJT_stage2_0.vr BGR_BJT_stage1_0.vr.t20 26.0492
R179 BGR_BJT_stage1_0.vr.n1 BGR_BJT_stage1_0.vr.n12 24.2089
R180 BGR_BJT_stage1_0.vr.n2 BGR_BJT_stage1_0.vr.n6 23.2516
R181 BGR_BJT_stage1_0.vr.n2 BGR_BJT_stage1_0.vr.n7 23.2516
R182 BGR_BJT_stage1_0.vr.n2 BGR_BJT_stage1_0.vr.n8 23.2516
R183 BGR_BJT_stage1_0.vr.n1 BGR_BJT_stage1_0.vr.n9 23.2516
R184 BGR_BJT_stage1_0.vr.n1 BGR_BJT_stage1_0.vr.n10 23.2516
R185 BGR_BJT_stage1_0.vr.n1 BGR_BJT_stage1_0.vr.n11 23.2516
R186 BGR_BJT_stage1_0.vr.n0 BGR_BJT_stage1_0.vr.t0 23
R187 BGR_BJT_stage1_0.vr.n0 BGR_BJT_stage1_0.vr.t2 23
R188 BGR_BJT_stage1_0.vr.n0 BGR_BJT_stage1_0.vr.n1 5.80801
R189 BGR_BJT_stage1_0.vr.n0 BGR_BJT_stage2_0.vr 4.90984
R190 BGR_BJT_stage1_0.vr.n1 BGR_BJT_stage1_0.vr.n2 4.51621
R191 BGR_BJT_stage1_0.vr.n6 BGR_BJT_stage1_0.vr.t18 4.3505
R192 BGR_BJT_stage1_0.vr.n6 BGR_BJT_stage1_0.vr.t11 4.3505
R193 BGR_BJT_stage1_0.vr.n7 BGR_BJT_stage1_0.vr.t6 4.3505
R194 BGR_BJT_stage1_0.vr.n7 BGR_BJT_stage1_0.vr.t14 4.3505
R195 BGR_BJT_stage1_0.vr.n8 BGR_BJT_stage1_0.vr.t15 4.3505
R196 BGR_BJT_stage1_0.vr.n8 BGR_BJT_stage1_0.vr.t12 4.3505
R197 BGR_BJT_stage1_0.vr.n9 BGR_BJT_stage1_0.vr.t13 4.3505
R198 BGR_BJT_stage1_0.vr.n9 BGR_BJT_stage1_0.vr.t10 4.3505
R199 BGR_BJT_stage1_0.vr.n10 BGR_BJT_stage1_0.vr.t16 4.3505
R200 BGR_BJT_stage1_0.vr.n10 BGR_BJT_stage1_0.vr.t7 4.3505
R201 BGR_BJT_stage1_0.vr.n11 BGR_BJT_stage1_0.vr.t9 4.3505
R202 BGR_BJT_stage1_0.vr.n11 BGR_BJT_stage1_0.vr.t5 4.3505
R203 BGR_BJT_stage1_0.vr.n12 BGR_BJT_stage1_0.vr.t4 4.3505
R204 BGR_BJT_stage1_0.vr.n12 BGR_BJT_stage1_0.vr.t17 4.3505
R205 BGR_BJT_stage1_0.vr.n4 BGR_BJT_stage1_0.vr.n3 2.80213
R206 BGR_BJT_stage2_0.vr BGR_BJT_stage1_0.vr.n5 2.76952
R207 BGR_BJT_stage1_0.vr.n5 BGR_BJT_stage1_0.vr.n4 2.72333
R208 BGR_BJT_stage1_0.vref0 BGR_BJT_stage1_0.vref0.t0 88.7532
R209 BGR_BJT_stage1_0.vref0.n16 BGR_BJT_stage1_0.vref0.n14 22.2005
R210 BGR_BJT_stage1_0.vref0.n6 BGR_BJT_stage1_0.vref0.n5 21.8815
R211 BGR_BJT_stage1_0.vref0.n6 BGR_BJT_stage1_0.vref0.n4 21.5624
R212 BGR_BJT_stage1_0.vref0.n9 BGR_BJT_stage1_0.vref0.n3 21.5624
R213 BGR_BJT_stage1_0.vref0.n10 BGR_BJT_stage1_0.vref0.n2 21.5624
R214 BGR_BJT_stage1_0.vref0.n11 BGR_BJT_stage1_0.vref0.n1 21.5624
R215 BGR_BJT_stage1_0.vref0.n0 BGR_BJT_stage1_0.vref0.n12 21.5624
R216 BGR_BJT_stage1_0.vref0.n8 BGR_BJT_stage1_0.vref0.n7 21.5624
R217 BGR_BJT_stage1_0.vref0.n29 BGR_BJT_stage1_0.vref0.n13 21.5603
R218 BGR_BJT_stage1_0.vref0.n28 BGR_BJT_stage1_0.vref0.n27 21.5445
R219 BGR_BJT_stage1_0.vref0.n26 BGR_BJT_stage1_0.vref0.n25 21.5445
R220 BGR_BJT_stage1_0.vref0.n24 BGR_BJT_stage1_0.vref0.n23 21.5445
R221 BGR_BJT_stage1_0.vref0.n22 BGR_BJT_stage1_0.vref0.n21 21.5445
R222 BGR_BJT_stage1_0.vref0.n20 BGR_BJT_stage1_0.vref0.n19 21.5445
R223 BGR_BJT_stage1_0.vref0.n18 BGR_BJT_stage1_0.vref0.n17 21.5445
R224 BGR_BJT_stage1_0.vref0.n16 BGR_BJT_stage1_0.vref0.n15 21.5445
R225 BGR_BJT_stage1_0.vref0.n5 BGR_BJT_stage1_0.vref0.t27 4.3505
R226 BGR_BJT_stage1_0.vref0.n5 BGR_BJT_stage1_0.vref0.t10 4.3505
R227 BGR_BJT_stage1_0.vref0.n4 BGR_BJT_stage1_0.vref0.t14 4.3505
R228 BGR_BJT_stage1_0.vref0.n4 BGR_BJT_stage1_0.vref0.t3 4.3505
R229 BGR_BJT_stage1_0.vref0.n3 BGR_BJT_stage1_0.vref0.t11 4.3505
R230 BGR_BJT_stage1_0.vref0.n3 BGR_BJT_stage1_0.vref0.t25 4.3505
R231 BGR_BJT_stage1_0.vref0.n2 BGR_BJT_stage1_0.vref0.t1 4.3505
R232 BGR_BJT_stage1_0.vref0.n2 BGR_BJT_stage1_0.vref0.t19 4.3505
R233 BGR_BJT_stage1_0.vref0.n1 BGR_BJT_stage1_0.vref0.t6 4.3505
R234 BGR_BJT_stage1_0.vref0.n1 BGR_BJT_stage1_0.vref0.t2 4.3505
R235 BGR_BJT_stage1_0.vref0.n12 BGR_BJT_stage1_0.vref0.t30 4.3505
R236 BGR_BJT_stage1_0.vref0.n12 BGR_BJT_stage1_0.vref0.t13 4.3505
R237 BGR_BJT_stage1_0.vref0.n13 BGR_BJT_stage1_0.vref0.t9 4.3505
R238 BGR_BJT_stage1_0.vref0.n13 BGR_BJT_stage1_0.vref0.t32 4.3505
R239 BGR_BJT_stage1_0.vref0.n27 BGR_BJT_stage1_0.vref0.t26 4.3505
R240 BGR_BJT_stage1_0.vref0.n27 BGR_BJT_stage1_0.vref0.t18 4.3505
R241 BGR_BJT_stage1_0.vref0.n25 BGR_BJT_stage1_0.vref0.t16 4.3505
R242 BGR_BJT_stage1_0.vref0.n25 BGR_BJT_stage1_0.vref0.t23 4.3505
R243 BGR_BJT_stage1_0.vref0.n23 BGR_BJT_stage1_0.vref0.t31 4.3505
R244 BGR_BJT_stage1_0.vref0.n23 BGR_BJT_stage1_0.vref0.t17 4.3505
R245 BGR_BJT_stage1_0.vref0.n21 BGR_BJT_stage1_0.vref0.t20 4.3505
R246 BGR_BJT_stage1_0.vref0.n21 BGR_BJT_stage1_0.vref0.t5 4.3505
R247 BGR_BJT_stage1_0.vref0.n19 BGR_BJT_stage1_0.vref0.t29 4.3505
R248 BGR_BJT_stage1_0.vref0.n19 BGR_BJT_stage1_0.vref0.t15 4.3505
R249 BGR_BJT_stage1_0.vref0.n17 BGR_BJT_stage1_0.vref0.t8 4.3505
R250 BGR_BJT_stage1_0.vref0.n17 BGR_BJT_stage1_0.vref0.t24 4.3505
R251 BGR_BJT_stage1_0.vref0.n15 BGR_BJT_stage1_0.vref0.t28 4.3505
R252 BGR_BJT_stage1_0.vref0.n15 BGR_BJT_stage1_0.vref0.t7 4.3505
R253 BGR_BJT_stage1_0.vref0.n14 BGR_BJT_stage1_0.vref0.t12 4.3505
R254 BGR_BJT_stage1_0.vref0.n14 BGR_BJT_stage1_0.vref0.t4 4.3505
R255 BGR_BJT_stage1_0.vref0.n7 BGR_BJT_stage1_0.vref0.t22 4.3505
R256 BGR_BJT_stage1_0.vref0.n7 BGR_BJT_stage1_0.vref0.t21 4.3505
R257 BGR_BJT_stage1_0.vref0.n29 BGR_BJT_stage1_0.vref0.n28 1.5282
R258 BGR_BJT_stage1_0.vref0.n8 BGR_BJT_stage1_0.vref0.n6 0.638711
R259 BGR_BJT_stage1_0.vref0.n10 BGR_BJT_stage1_0.vref0.n9 0.638711
R260 BGR_BJT_stage1_0.vref0.n20 BGR_BJT_stage1_0.vref0.n18 0.624699
R261 BGR_BJT_stage1_0.vref0.n24 BGR_BJT_stage1_0.vref0.n22 0.624699
R262 BGR_BJT_stage1_0.vref0.n28 BGR_BJT_stage1_0.vref0.n26 0.624699
R263 BGR_BJT_stage1_0.vref0.n0 BGR_BJT_stage1_0.vref0.n11 0.59171
R264 BGR_BJT_stage1_0.vref0 BGR_BJT_stage1_0.vref0.n0 0.435868
R265 BGR_BJT_stage1_0.vref0.n0 BGR_BJT_stage1_0.vref0.n29 0.366605
R266 BGR_BJT_stage1_0.vref0.n9 BGR_BJT_stage1_0.vref0.n8 0.319605
R267 BGR_BJT_stage1_0.vref0.n11 BGR_BJT_stage1_0.vref0.n10 0.319605
R268 BGR_BJT_stage1_0.vref0.n18 BGR_BJT_stage1_0.vref0.n16 0.296969
R269 BGR_BJT_stage1_0.vref0.n22 BGR_BJT_stage1_0.vref0.n20 0.296969
R270 BGR_BJT_stage1_0.vref0.n26 BGR_BJT_stage1_0.vref0.n24 0.296969
R271 vss.t43 vss.n38 310750
R272 vss.n262 vss.n38 224782
R273 vss.n268 vss.n264 133392
R274 vss.n262 vss.n261 52883
R275 vss.n20 vss.n19 26954.2
R276 vss.n277 vss.n19 26954.2
R277 vss.n276 vss.n20 26948.4
R278 vss.n277 vss.n276 26948.4
R279 vss.n269 vss.n23 17753.2
R280 vss.n273 vss.n23 17753.2
R281 vss.n273 vss.n24 17753.2
R282 vss.n269 vss.n24 17753.2
R283 vss.n263 vss.n262 11463.8
R284 vss.n264 vss.n263 9418.38
R285 vss.n177 vss.n17 7283.2
R286 vss.n263 vss.n22 7271.49
R287 vss.n265 vss.n264 7271.49
R288 vss.n177 vss.n44 6748.27
R289 vss.n107 vss.n25 3062.16
R290 vss.n261 vss.n39 1611.76
R291 vss.n231 vss.n64 1517.24
R292 vss.n221 vss.n64 1517.24
R293 vss.n221 vss.n59 1517.24
R294 vss.n233 vss.n59 1517.24
R295 vss.n246 vss.n51 1517.24
R296 vss.n247 vss.n246 1517.24
R297 vss.n248 vss.n247 1517.24
R298 vss.n248 vss.n40 1517.24
R299 vss.n260 vss.n40 1517.24
R300 vss.n232 vss.n231 1489.48
R301 vss.n89 vss.n18 1058.82
R302 vss.n170 vss.n89 1058.82
R303 vss.n171 vss.n170 1058.82
R304 vss.n172 vss.n171 1058.82
R305 vss.n172 vss.n60 1058.82
R306 vss.n193 vss.n61 1058.82
R307 vss.n193 vss.n192 1058.82
R308 vss.n192 vss.n191 1058.82
R309 vss.n191 vss.n187 1058.82
R310 vss.n187 vss.n39 1058.82
R311 vss.t43 vss.n51 792.337
R312 vss.n233 vss.t43 724.904
R313 vss.t43 vss.n61 717.648
R314 vss.n232 vss.n63 599.813
R315 vss.n278 vss.n18 591.216
R316 vss.n280 vss.n14 585
R317 vss.n283 vss.n282 585
R318 vss.n279 vss.n17 585
R319 vss.n279 vss.n278 585
R320 vss.n91 vss.n16 585
R321 vss.n18 vss.n16 585
R322 vss.n156 vss.n12 585
R323 vss.n284 vss.n12 585
R324 vss.n287 vss.n286 585
R325 vss.n286 vss.n285 585
R326 vss.n150 vss.n11 585
R327 vss.n13 vss.n11 585
R328 vss.n149 vss.n148 585
R329 vss.n148 vss.n147 585
R330 vss.n101 vss.n97 585
R331 vss.n146 vss.n97 585
R332 vss.n144 vss.n143 585
R333 vss.n145 vss.n144 585
R334 vss.n135 vss.n99 585
R335 vss.n99 vss.n98 585
R336 vss.n134 vss.n133 585
R337 vss.n133 vss.n132 585
R338 vss.n127 vss.n104 585
R339 vss.n131 vss.n104 585
R340 vss.n129 vss.n128 585
R341 vss.n130 vss.n129 585
R342 vss.n107 vss.n106 585
R343 vss.n106 vss.n62 585
R344 vss.n122 vss.n107 585
R345 vss.n125 vss.n124 585
R346 vss.n121 vss.n120 585
R347 vss.n114 vss.n113 585
R348 vss.n112 vss.n81 585
R349 vss.n200 vss.n78 585
R350 vss.n209 vss.n208 585
R351 vss.n211 vss.n77 585
R352 vss.n212 vss.n70 585
R353 vss.n215 vss.n214 585
R354 vss.n75 vss.n74 585
R355 vss.n74 vss.n73 585
R356 vss.n42 vss.n39 585
R357 vss.n189 vss.n187 585
R358 vss.n259 vss.n258 585
R359 vss.n260 vss.n259 585
R360 vss.n43 vss.n41 585
R361 vss.n41 vss.n40 585
R362 vss.n250 vss.n249 585
R363 vss.n249 vss.n248 585
R364 vss.n50 vss.n49 585
R365 vss.n247 vss.n50 585
R366 vss.n245 vss.n244 585
R367 vss.n246 vss.n245 585
R368 vss.n54 vss.n52 585
R369 vss.n52 vss.n51 585
R370 vss.n235 vss.n234 585
R371 vss.n234 vss.n233 585
R372 vss.n58 vss.n57 585
R373 vss.n59 vss.n58 585
R374 vss.n223 vss.n222 585
R375 vss.n222 vss.n221 585
R376 vss.n67 vss.n65 585
R377 vss.n65 vss.n64 585
R378 vss.n230 vss.n229 585
R379 vss.n231 vss.n230 585
R380 vss.n66 vss.n63 585
R381 vss.n190 vss.n45 585
R382 vss.n191 vss.n190 585
R383 vss.n186 vss.n185 585
R384 vss.n192 vss.n186 585
R385 vss.n195 vss.n194 585
R386 vss.n194 vss.n193 585
R387 vss.n176 vss.n84 585
R388 vss.n84 vss.n61 585
R389 vss.n175 vss.n174 585
R390 vss.n174 vss.n60 585
R391 vss.n173 vss.n88 585
R392 vss.n173 vss.n172 585
R393 vss.n94 vss.n87 585
R394 vss.n171 vss.n87 585
R395 vss.n169 vss.n168 585
R396 vss.n170 vss.n169 585
R397 vss.n92 vss.n90 585
R398 vss.n90 vss.n89 585
R399 vss.t43 vss.n232 369.531
R400 vss.n269 vss.t41 343.529
R401 vss.t43 vss.n60 341.176
R402 vss.n261 vss.n260 337.166
R403 vss.n272 vss.n271 281.336
R404 vss.n271 vss.n270 281.243
R405 vss.n255 vss.n254 258.334
R406 vss.n73 vss.n63 257.466
R407 vss.n26 vss.n6 255.369
R408 vss.n281 vss.n15 254.34
R409 vss.n123 vss.n62 254.34
R410 vss.n109 vss.n62 254.34
R411 vss.n111 vss.n62 254.34
R412 vss.n210 vss.n62 254.34
R413 vss.n213 vss.n62 254.34
R414 vss.n71 vss.n62 254.34
R415 vss.n188 vss.n44 254.34
R416 vss.n259 vss.n42 251.614
R417 vss.n227 vss.n219 250
R418 vss.t41 vss.t37 242.773
R419 vss.t37 vss.t39 242.773
R420 vss.t52 vss.t21 242.773
R421 vss.t50 vss.n274 203.251
R422 vss.n157 vss.n7 200.249
R423 vss.n38 vss.t23 195.724
R424 vss.n129 vss.n105 195.049
R425 vss.n280 vss.n279 187.249
R426 vss.n159 vss.n158 185
R427 vss.n155 vss.n10 185
R428 vss.n155 vss.t42 185
R429 vss.n154 vss.n9 185
R430 vss.n152 vss.n151 185
R431 vss.n96 vss.n95 185
R432 vss.n142 vss.n141 185
R433 vss.n139 vss.n100 185
R434 vss.n137 vss.n136 185
R435 vss.n103 vss.n102 185
R436 vss.n116 vss.n108 185
R437 vss.n119 vss.n118 185
R438 vss.n110 vss.n80 185
R439 vss.n202 vss.n201 185
R440 vss.n204 vss.n79 185
R441 vss.n207 vss.n206 185
R442 vss.n76 vss.n69 185
R443 vss.n217 vss.n216 185
R444 vss.n219 vss.n68 185
R445 vss.n254 vss.n47 185
R446 vss.n252 vss.n251 185
R447 vss.n243 vss.n48 185
R448 vss.n242 vss.n241 185
R449 vss.n239 vss.n55 185
R450 vss.n237 vss.n236 185
R451 vss.n220 vss.n56 185
R452 vss.n56 vss.t42 185
R453 vss.n225 vss.n224 185
R454 vss.n228 vss.n227 185
R455 vss.n256 vss.n255 185
R456 vss.n184 vss.n183 185
R457 vss.n182 vss.n83 185
R458 vss.n180 vss.n82 185
R459 vss.n179 vss.n178 185
R460 vss.n162 vss.n86 185
R461 vss.n164 vss.n163 185
R462 vss.n167 vss.n166 185
R463 vss.n161 vss.n93 185
R464 vss.n267 vss.t40 181.608
R465 vss.n90 vss.n16 175.546
R466 vss.n169 vss.n90 175.546
R467 vss.n169 vss.n87 175.546
R468 vss.n173 vss.n87 175.546
R469 vss.n174 vss.n173 175.546
R470 vss.n174 vss.n84 175.546
R471 vss.n194 vss.n84 175.546
R472 vss.n194 vss.n186 175.546
R473 vss.n190 vss.n186 175.546
R474 vss.n190 vss.n189 175.546
R475 vss.n230 vss.n63 175.546
R476 vss.n230 vss.n65 175.546
R477 vss.n222 vss.n65 175.546
R478 vss.n222 vss.n58 175.546
R479 vss.n234 vss.n58 175.546
R480 vss.n234 vss.n52 175.546
R481 vss.n245 vss.n52 175.546
R482 vss.n245 vss.n50 175.546
R483 vss.n249 vss.n50 175.546
R484 vss.n249 vss.n41 175.546
R485 vss.n259 vss.n41 175.546
R486 vss.n124 vss.n121 175.546
R487 vss.n113 vss.n112 175.546
R488 vss.n209 vss.n78 175.546
R489 vss.n212 vss.n211 175.546
R490 vss.n214 vss.n75 175.546
R491 vss.n129 vss.n104 175.546
R492 vss.n133 vss.n104 175.546
R493 vss.n133 vss.n99 175.546
R494 vss.n144 vss.n99 175.546
R495 vss.n144 vss.n97 175.546
R496 vss.n148 vss.n97 175.546
R497 vss.n148 vss.n11 175.546
R498 vss.n286 vss.n11 175.546
R499 vss.n286 vss.n12 175.546
R500 vss.n282 vss.n12 175.546
R501 vss.n62 vss.t52 169.376
R502 vss.t25 vss.t38 167.494
R503 vss.t53 vss.t57 167.494
R504 vss.t19 vss.t59 167.494
R505 vss.t27 vss.t60 167.494
R506 vss.t54 vss.t58 167.494
R507 vss.t0 vss.t56 167.494
R508 vss.t49 vss.t13 167.494
R509 vss.t8 vss.t12 167.494
R510 vss.t29 vss.t15 167.494
R511 vss.t55 vss.t14 167.494
R512 vss.t6 vss.t47 167.494
R513 vss.t51 vss.t44 167.494
R514 vss.t10 vss.t45 167.494
R515 vss.t2 vss.t48 167.494
R516 vss.n166 vss.n161 150
R517 vss.n164 vss.n162 150
R518 vss.n180 vss.n179 150
R519 vss.n183 vss.n182 150
R520 vss.n225 vss.n56 150
R521 vss.n237 vss.n56 150
R522 vss.n241 vss.n239 150
R523 vss.n252 vss.n48 150
R524 vss.n118 vss.n116 150
R525 vss.n202 vss.n80 150
R526 vss.n206 vss.n204 150
R527 vss.n217 vss.n69 150
R528 vss.n137 vss.n102 150
R529 vss.n141 vss.n139 150
R530 vss.n152 vss.n95 150
R531 vss.n155 vss.n154 150
R532 vss.n159 vss.n155 150
R533 vss.n37 vss.n26 147.531
R534 vss.t31 vss.n22 140.206
R535 vss.n293 vss.n292 137.462
R536 vss.n279 vss.n16 126.782
R537 vss.n122 vss.n105 124.832
R538 vss.n278 vss.n14 124.675
R539 vss.n294 vss.n293 122.373
R540 vss.n131 vss.n130 116.883
R541 vss.n132 vss.n131 116.883
R542 vss.n145 vss.n98 116.883
R543 vss.n146 vss.n145 116.883
R544 vss.n147 vss.n13 116.883
R545 vss.n285 vss.n13 116.883
R546 vss.n284 vss.n283 116.883
R547 vss.n283 vss.n14 116.883
R548 vss.n266 vss.n265 94.098
R549 vss.t35 vss.n284 76.6239
R550 vss.n188 vss.n42 76.3222
R551 vss.n123 vss.n122 76.3222
R552 vss.n121 vss.n109 76.3222
R553 vss.n112 vss.n111 76.3222
R554 vss.n210 vss.n209 76.3222
R555 vss.n213 vss.n212 76.3222
R556 vss.n75 vss.n71 76.3222
R557 vss.n281 vss.n280 76.3222
R558 vss.n282 vss.n281 76.3222
R559 vss.n124 vss.n123 76.3222
R560 vss.n113 vss.n109 76.3222
R561 vss.n111 vss.n78 76.3222
R562 vss.n211 vss.n210 76.3222
R563 vss.n214 vss.n213 76.3222
R564 vss.n73 vss.n71 76.3222
R565 vss.n189 vss.n188 76.3222
R566 vss.t40 vss.t25 75.2785
R567 vss.t38 vss.t53 75.2785
R568 vss.t57 vss.t19 75.2785
R569 vss.t59 vss.t27 75.2785
R570 vss.t60 vss.t54 75.2785
R571 vss.t58 vss.t0 75.2785
R572 vss.t56 vss.t17 75.2785
R573 vss.t16 vss.t49 75.2785
R574 vss.t13 vss.t8 75.2785
R575 vss.t12 vss.t29 75.2785
R576 vss.t15 vss.t55 75.2785
R577 vss.t14 vss.t31 75.2785
R578 vss.t46 vss.t6 75.2785
R579 vss.t47 vss.t51 75.2785
R580 vss.t44 vss.t10 75.2785
R581 vss.t45 vss.t2 75.2785
R582 vss.t48 vss.t50 75.2785
R583 vss.t43 vss.n62 72.4556
R584 vss.n132 vss.t4 71.4291
R585 vss.n161 vss.n160 69.3109
R586 vss.n160 vss.n159 69.3109
R587 vss.n270 vss.n37 66.0923
R588 vss.n153 vss.t42 65.8183
R589 vss.n140 vss.t42 65.8183
R590 vss.n138 vss.t42 65.8183
R591 vss.n117 vss.t42 65.8183
R592 vss.n203 vss.t42 65.8183
R593 vss.n205 vss.t42 65.8183
R594 vss.n218 vss.t42 65.8183
R595 vss.n253 vss.t42 65.8183
R596 vss.n240 vss.t42 65.8183
R597 vss.n238 vss.t42 65.8183
R598 vss.n226 vss.t42 65.8183
R599 vss.t42 vss.n46 65.8183
R600 vss.n181 vss.t42 65.8183
R601 vss.n85 vss.t42 65.8183
R602 vss.n165 vss.t42 65.8183
R603 vss.n270 vss.n269 65.0005
R604 vss.n273 vss.n272 65.0005
R605 vss.n274 vss.n273 65.0005
R606 vss.n115 vss.t42 64.1729
R607 vss.n147 vss.t43 61.0395
R608 vss.n160 vss.t42 57.8461
R609 vss.n116 vss.n115 56.6572
R610 vss.n115 vss.n102 56.6572
R611 vss.t43 vss.n146 55.8447
R612 vss.n165 vss.n164 53.3664
R613 vss.n179 vss.n85 53.3664
R614 vss.n182 vss.n181 53.3664
R615 vss.n255 vss.n46 53.3664
R616 vss.n227 vss.n226 53.3664
R617 vss.n238 vss.n237 53.3664
R618 vss.n241 vss.n240 53.3664
R619 vss.n253 vss.n252 53.3664
R620 vss.n118 vss.n117 53.3664
R621 vss.n203 vss.n202 53.3664
R622 vss.n206 vss.n205 53.3664
R623 vss.n218 vss.n217 53.3664
R624 vss.n138 vss.n137 53.3664
R625 vss.n141 vss.n140 53.3664
R626 vss.n153 vss.n152 53.3664
R627 vss.n154 vss.n153 53.3664
R628 vss.n140 vss.n95 53.3664
R629 vss.n139 vss.n138 53.3664
R630 vss.n117 vss.n80 53.3664
R631 vss.n204 vss.n203 53.3664
R632 vss.n205 vss.n69 53.3664
R633 vss.n219 vss.n218 53.3664
R634 vss.n254 vss.n253 53.3664
R635 vss.n240 vss.n48 53.3664
R636 vss.n239 vss.n238 53.3664
R637 vss.n226 vss.n225 53.3664
R638 vss.n183 vss.n46 53.3664
R639 vss.n181 vss.n180 53.3664
R640 vss.n162 vss.n85 53.3664
R641 vss.n166 vss.n165 53.3664
R642 vss.n268 vss.n267 52.6951
R643 vss.t21 vss.n38 47.0493
R644 vss.t17 vss.n266 46.1083
R645 vss.t4 vss.n98 45.455
R646 vss.n285 vss.t35 40.2602
R647 vss.n274 vss.t23 39.5215
R648 vss.n292 vss.n7 32.2788
R649 vss.n130 vss.t33 29.8706
R650 vss.n265 vss.t16 27.2888
R651 vss.n28 vss.t26 26.5035
R652 vss.n290 vss.t36 25.0376
R653 vss.n272 vss.n25 23.4151
R654 vss.n37 vss.n36 23.2185
R655 vss.n5 vss.n4 21.6664
R656 vss.n28 vss.n27 20.6876
R657 vss.n32 vss.n29 20.6876
R658 vss.n31 vss.n30 20.6876
R659 vss.n297 vss.n1 20.6683
R660 vss.n296 vss.n2 20.6683
R661 vss.n5 vss.n3 20.6683
R662 vss.n275 vss.t46 16.9381
R663 vss.n25 vss.n21 16.9125
R664 vss.n35 vss.n34 16.6367
R665 vss.n277 vss.n7 14.6255
R666 vss.n278 vss.n277 14.6255
R667 vss.n26 vss.n20 14.6255
R668 vss.n267 vss.n20 14.6255
R669 vss.n275 vss.n22 10.3512
R670 vss.t39 vss.n268 8.46928
R671 vss.n271 vss.n24 7.313
R672 vss.n266 vss.n24 7.313
R673 vss.n36 vss.n23 7.313
R674 vss.n266 vss.n23 7.313
R675 vss.n292 vss.n291 6.9005
R676 vss.n293 vss.n0 6.9005
R677 vss.n19 vss.n6 6.15839
R678 vss.n275 vss.n19 6.15839
R679 vss.n276 vss.n21 6.15839
R680 vss.n276 vss.n275 6.15839
R681 vss.n229 vss.n66 4.90263
R682 vss.n258 vss.n43 4.90263
R683 vss.n168 vss.n93 4.88977
R684 vss.n167 vss.n94 4.88977
R685 vss.n163 vss.n88 4.88977
R686 vss.n175 vss.n86 4.88977
R687 vss.n185 vss.n83 4.88977
R688 vss.n184 vss.n45 4.88977
R689 vss.n92 vss.n91 4.65477
R690 vss.n91 vss.n17 4.57193
R691 vss.n27 vss.t1 4.3505
R692 vss.n27 vss.t18 4.3505
R693 vss.n29 vss.t32 4.3505
R694 vss.n29 vss.t7 4.3505
R695 vss.n30 vss.t24 4.3505
R696 vss.n30 vss.t22 4.3505
R697 vss.n1 vss.t34 4.3505
R698 vss.n1 vss.t5 4.3505
R699 vss.n2 vss.t11 4.3505
R700 vss.n2 vss.t3 4.3505
R701 vss.n3 vss.t9 4.3505
R702 vss.n3 vss.t30 4.3505
R703 vss.n4 vss.t20 4.3505
R704 vss.n4 vss.t28 4.3505
R705 vss.n257 vss.n256 4.23054
R706 vss.n291 vss.n290 4.10351
R707 vss.n157 vss.n15 3.9624
R708 vss.n120 vss.n108 3.81327
R709 vss.n119 vss.n114 3.81327
R710 vss.n110 vss.n81 3.81327
R711 vss.n201 vss.n200 3.81327
R712 vss.n208 vss.n79 3.81327
R713 vss.n207 vss.n77 3.81327
R714 vss.n76 vss.n70 3.81327
R715 vss.n216 vss.n215 3.81327
R716 vss.n74 vss.n72 3.70433
R717 vss.n257 vss.n44 3.64986
R718 vss.n196 vss.n82 3.57132
R719 vss.n177 vss.n176 3.35157
R720 vss.n72 vss.n68 3.15965
R721 vss.n229 vss.n228 2.7239
R722 vss.n224 vss.n67 2.7239
R723 vss.n223 vss.n220 2.7239
R724 vss.n236 vss.n57 2.7239
R725 vss.n235 vss.n55 2.7239
R726 vss.n244 vss.n243 2.7239
R727 vss.n251 vss.n49 2.7239
R728 vss.n250 vss.n47 2.7239
R729 vss.n291 vss.n0 2.28754
R730 vss.n228 vss.n67 2.17922
R731 vss.n224 vss.n223 2.17922
R732 vss.n220 vss.n57 2.17922
R733 vss.n236 vss.n235 2.17922
R734 vss.n55 vss.n54 2.17922
R735 vss.n244 vss.n242 2.17922
R736 vss.n243 vss.n49 2.17922
R737 vss.n251 vss.n250 2.17922
R738 vss.n47 vss.n43 2.17922
R739 vss.n128 vss.n127 2.17819
R740 vss.n106 vss.n105 1.951
R741 vss.n289 vss.n288 1.89157
R742 vss.n72 vss.n66 1.79795
R743 vss.n134 vss.n103 1.79105
R744 vss.n136 vss.n135 1.79105
R745 vss.n143 vss.n100 1.79105
R746 vss.n142 vss.n101 1.79105
R747 vss.n149 vss.n96 1.79105
R748 vss.n156 vss.n10 1.79105
R749 vss.n35 vss 1.7155
R750 vss.n54 vss.n53 1.68901
R751 vss.n126 vss.n107 1.64587
R752 vss.n258 vss.n257 1.58007
R753 vss.n178 vss.n177 1.5387
R754 vss.n197 vss.n196 1.519
R755 vss.n32 vss.n31 1.46641
R756 vss.n33 vss.n28 1.43989
R757 vss vss.n150 1.37971
R758 vss.n158 vss.n157 1.37971
R759 vss.n196 vss.n195 1.31895
R760 vss.n288 vss.n287 1.18613
R761 vss.n17 vss.n15 1.16875
R762 vss.n126 vss.n125 1.08986
R763 vss.n125 vss.n108 1.08986
R764 vss.n120 vss.n119 1.08986
R765 vss.n114 vss.n110 1.08986
R766 vss.n201 vss.n81 1.08986
R767 vss.n208 vss.n207 1.08986
R768 vss.n77 vss.n76 1.08986
R769 vss.n216 vss.n70 1.08986
R770 vss.n215 vss.n68 1.08986
R771 vss.n242 vss.n53 1.03539
R772 vss.n297 vss.n296 0.997923
R773 vss.n199 vss.n79 0.817521
R774 vss.n128 vss.n126 0.798988
R775 vss.n198 vss.n197 0.76482
R776 vss.n34 vss.n21 0.740167
R777 vss.n198 vss.n8 0.654721
R778 vss.n298 vss.n297 0.633876
R779 vss.n288 vss.n9 0.605415
R780 vss.n197 vss.n53 0.596304
R781 vss.n199 vss.n198 0.59175
R782 vss.t43 vss.t33 0.546135
R783 vss.n31 vss.n8 0.539326
R784 vss.n294 vss.n6 0.532356
R785 vss.n295 vss.n5 0.528206
R786 vss.n296 vss.n295 0.469572
R787 vss.n289 vss.n8 0.452967
R788 vss.n151 vss 0.411842
R789 vss.n127 vss.n103 0.387646
R790 vss.n136 vss.n134 0.387646
R791 vss.n135 vss.n100 0.387646
R792 vss.n143 vss.n142 0.387646
R793 vss.n101 vss.n96 0.387646
R794 vss.n150 vss.n9 0.387646
R795 vss.n287 vss.n10 0.387646
R796 vss.n158 vss.n156 0.387646
R797 vss.n298 vss.n0 0.343093
R798 vss.n200 vss.n199 0.27284
R799 vss vss.n149 0.242466
R800 vss.n36 vss.n35 0.188551
R801 vss.n151 vss 0.14568
R802 vss.n34 vss.n33 0.0987955
R803 vss.n290 vss.n289 0.0948141
R804 vss vss.n298 0.0849072
R805 vss.n295 vss.n294 0.0736577
R806 vss.n93 vss.n92 0.0554356
R807 vss.n168 vss.n167 0.0554356
R808 vss.n163 vss.n94 0.0554356
R809 vss.n88 vss.n86 0.0554356
R810 vss.n178 vss.n175 0.0554356
R811 vss.n176 vss.n82 0.0554356
R812 vss.n195 vss.n83 0.0554356
R813 vss.n185 vss.n184 0.0554356
R814 vss.n256 vss.n45 0.0554356
R815 vss.n33 vss.n32 0.0270152
R816 a_365_2822.n24 a_365_2822.t18 190.305
R817 a_365_2822.t18 a_365_2822.n23 190.305
R818 a_365_2822.n25 a_365_2822.t26 190.305
R819 a_365_2822.t26 a_365_2822.n21 190.305
R820 a_365_2822.n42 a_365_2822.t28 190.305
R821 a_365_2822.n34 a_365_2822.t28 190.305
R822 a_365_2822.n38 a_365_2822.t16 190.305
R823 a_365_2822.t16 a_365_2822.n33 190.305
R824 a_365_2822.n62 a_365_2822.t4 190.305
R825 a_365_2822.t4 a_365_2822.n44 190.305
R826 a_365_2822.t6 a_365_2822.n63 190.305
R827 a_365_2822.n64 a_365_2822.t6 190.305
R828 a_365_2822.n67 a_365_2822.t0 190.305
R829 a_365_2822.t0 a_365_2822.n29 190.305
R830 a_365_2822.n32 a_365_2822.t10 190.305
R831 a_365_2822.t10 a_365_2822.n31 190.305
R832 a_365_2822.n50 a_365_2822.t2 190.305
R833 a_365_2822.t2 a_365_2822.n15 190.305
R834 a_365_2822.n51 a_365_2822.t14 190.305
R835 a_365_2822.t14 a_365_2822.n14 190.305
R836 a_365_2822.n74 a_365_2822.t8 190.305
R837 a_365_2822.n19 a_365_2822.t8 190.305
R838 a_365_2822.t20 a_365_2822.n18 190.305
R839 a_365_2822.n71 a_365_2822.t20 190.305
R840 a_365_2822.n80 a_365_2822.t24 190.305
R841 a_365_2822.t24 a_365_2822.n79 190.305
R842 a_365_2822.n81 a_365_2822.t22 190.305
R843 a_365_2822.t22 a_365_2822.n77 190.305
R844 a_365_2822.n16 a_365_2822.t30 95.1811
R845 a_365_2822.n57 a_365_2822.t12 95.1783
R846 a_365_2822.n40 a_365_2822.n37 22.3176
R847 a_365_2822.n48 a_365_2822.n47 22.2301
R848 a_365_2822.n59 a_365_2822.n58 22.2284
R849 a_365_2822.n10 a_365_2822.n60 22.2284
R850 a_365_2822.n55 a_365_2822.n54 22.2284
R851 a_365_2822.n11 a_365_2822.n53 22.2284
R852 a_365_2822.n7 a_365_2822.n46 22.2284
R853 a_365_2822.n1 a_365_2822.n83 22.2284
R854 a_365_2822.n84 a_365_2822.n4 22.2284
R855 a_365_2822.n6 a_365_2822.n36 22.1884
R856 a_365_2822.n9 a_365_2822.n35 22.1884
R857 a_365_2822.n2 a_365_2822.n69 22.1884
R858 a_365_2822.n3 a_365_2822.n70 22.1884
R859 a_365_2822.n0 a_365_2822.n28 22.1884
R860 a_365_2822.n8 a_365_2822.n27 22.1884
R861 a_365_2822.n5 a_365_2822.n20 22.1884
R862 a_365_2822.n57 a_365_2822.n43 11.5566
R863 a_365_2822.n17 a_365_2822.n16 10.9335
R864 a_365_2822.n43 a_365_2822.n42 9.80925
R865 a_365_2822.n67 a_365_2822.n66 9.80925
R866 a_365_2822.n75 a_365_2822.n74 9.80925
R867 a_365_2822.n24 a_365_2822.n17 9.80925
R868 a_365_2822.n15 a_365_2822.n12 9.403
R869 a_365_2822.n65 a_365_2822.n64 9.39819
R870 a_365_2822.n77 a_365_2822.n76 9.39819
R871 a_365_2822.n59 a_365_2822.n57 4.9275
R872 a_365_2822.n16 a_365_2822.n4 4.79654
R873 a_365_2822.n22 a_365_2822.n5 4.5005
R874 a_365_2822.n8 a_365_2822.n26 4.5005
R875 a_365_2822.n73 a_365_2822.n0 4.5005
R876 a_365_2822.n3 a_365_2822.n72 4.5005
R877 a_365_2822.n2 a_365_2822.n68 4.5005
R878 a_365_2822.n30 a_365_2822.n9 4.5005
R879 a_365_2822.n41 a_365_2822.n6 4.5005
R880 a_365_2822.n40 a_365_2822.n39 4.5005
R881 a_365_2822.n1 a_365_2822.n82 4.5005
R882 a_365_2822.n78 a_365_2822.n7 4.5005
R883 a_365_2822.n13 a_365_2822.n49 4.5005
R884 a_365_2822.n11 a_365_2822.n52 4.5005
R885 a_365_2822.n56 a_365_2822.n45 4.5005
R886 a_365_2822.n61 a_365_2822.n10 4.5005
R887 a_365_2822.n58 a_365_2822.t37 4.3505
R888 a_365_2822.n58 a_365_2822.t13 4.3505
R889 a_365_2822.n60 a_365_2822.t5 4.3505
R890 a_365_2822.n60 a_365_2822.t35 4.3505
R891 a_365_2822.n54 a_365_2822.t41 4.3505
R892 a_365_2822.n54 a_365_2822.t7 4.3505
R893 a_365_2822.n53 a_365_2822.t15 4.3505
R894 a_365_2822.n53 a_365_2822.t44 4.3505
R895 a_365_2822.n47 a_365_2822.t39 4.3505
R896 a_365_2822.n47 a_365_2822.t3 4.3505
R897 a_365_2822.n46 a_365_2822.t25 4.3505
R898 a_365_2822.n46 a_365_2822.t43 4.3505
R899 a_365_2822.n83 a_365_2822.t38 4.3505
R900 a_365_2822.n83 a_365_2822.t23 4.3505
R901 a_365_2822.n37 a_365_2822.t17 4.3505
R902 a_365_2822.n37 a_365_2822.t42 4.3505
R903 a_365_2822.n36 a_365_2822.t40 4.3505
R904 a_365_2822.n36 a_365_2822.t29 4.3505
R905 a_365_2822.n35 a_365_2822.t11 4.3505
R906 a_365_2822.n35 a_365_2822.t33 4.3505
R907 a_365_2822.n69 a_365_2822.t34 4.3505
R908 a_365_2822.n69 a_365_2822.t1 4.3505
R909 a_365_2822.n70 a_365_2822.t21 4.3505
R910 a_365_2822.n70 a_365_2822.t46 4.3505
R911 a_365_2822.n28 a_365_2822.t32 4.3505
R912 a_365_2822.n28 a_365_2822.t9 4.3505
R913 a_365_2822.n27 a_365_2822.t27 4.3505
R914 a_365_2822.n27 a_365_2822.t45 4.3505
R915 a_365_2822.n20 a_365_2822.t36 4.3505
R916 a_365_2822.n20 a_365_2822.t19 4.3505
R917 a_365_2822.t31 a_365_2822.n84 4.3505
R918 a_365_2822.n84 a_365_2822.t47 4.3505
R919 a_365_2822.n5 a_365_2822.n4 2.55258
R920 a_365_2822.n76 a_365_2822.n17 1.86108
R921 a_365_2822.n76 a_365_2822.n75 1.86108
R922 a_365_2822.n75 a_365_2822.n12 1.86108
R923 a_365_2822.n66 a_365_2822.n12 1.86108
R924 a_365_2822.n66 a_365_2822.n65 1.86108
R925 a_365_2822.n65 a_365_2822.n43 1.86108
R926 a_365_2822.n4 a_365_2822.n1 1.20675
R927 a_365_2822.n0 a_365_2822.n8 1.0755
R928 a_365_2822.n3 a_365_2822.n2 1.0755
R929 a_365_2822.n6 a_365_2822.n9 1.0755
R930 a_365_2822.n48 a_365_2822.n7 1.0755
R931 a_365_2822.n55 a_365_2822.n11 1.0755
R932 a_365_2822.n10 a_365_2822.n59 1.0755
R933 a_365_2822.n52 a_365_2822.n51 0.759759
R934 a_365_2822.n50 a_365_2822.n13 0.756673
R935 a_365_2822.n63 a_365_2822.n45 0.702205
R936 a_365_2822.n62 a_365_2822.n61 0.700784
R937 a_365_2822.n72 a_365_2822.n71 0.669534
R938 a_365_2822.n68 a_365_2822.n29 0.668114
R939 a_365_2822.n41 a_365_2822.n34 0.666693
R940 a_365_2822.n73 a_365_2822.n19 0.665273
R941 a_365_2822.n26 a_365_2822.n21 0.662432
R942 a_365_2822.n23 a_365_2822.n22 0.662432
R943 a_365_2822.n39 a_365_2822.n38 0.659208
R944 a_365_2822.n52 a_365_2822.n14 0.645562
R945 a_365_2822.n15 a_365_2822.n13 0.645562
R946 a_365_2822.n26 a_365_2822.n25 0.631182
R947 a_365_2822.n24 a_365_2822.n22 0.631181
R948 a_365_2822.n31 a_365_2822.n30 0.629532
R949 a_365_2822.n74 a_365_2822.n73 0.62834
R950 a_365_2822.n42 a_365_2822.n41 0.626919
R951 a_365_2822.n68 a_365_2822.n67 0.625499
R952 a_365_2822.n72 a_365_2822.n18 0.62408
R953 a_365_2822.n39 a_365_2822.n33 0.619882
R954 a_365_2822.n32 a_365_2822.n30 0.594586
R955 a_365_2822.n61 a_365_2822.n44 0.59283
R956 a_365_2822.n64 a_365_2822.n45 0.591403
R957 a_365_2822.n82 a_365_2822.n81 0.580689
R958 a_365_2822.n80 a_365_2822.n78 0.57833
R959 a_365_2822.n8 a_365_2822.n5 0.538
R960 a_365_2822.n2 a_365_2822.n9 0.538
R961 a_365_2822.n1 a_365_2822.n7 0.538
R962 a_365_2822.n0 a_365_2822.n3 0.538
R963 a_365_2822.n79 a_365_2822.n78 0.495783
R964 a_365_2822.n82 a_365_2822.n77 0.493421
R965 a_365_2822.n15 a_365_2822.n14 0.490992
R966 a_365_2822.n51 a_365_2822.n50 0.486913
R967 a_365_2822.n42 a_365_2822.n33 0.476043
R968 a_365_2822.n38 a_365_2822.n34 0.476043
R969 a_365_2822.n25 a_365_2822.n24 0.459739
R970 a_365_2822.n23 a_365_2822.n21 0.459739
R971 a_365_2822.n67 a_365_2822.n32 0.459739
R972 a_365_2822.n31 a_365_2822.n29 0.459739
R973 a_365_2822.n74 a_365_2822.n18 0.459739
R974 a_365_2822.n71 a_365_2822.n19 0.459739
R975 a_365_2822.n64 a_365_2822.n44 0.451587
R976 a_365_2822.n63 a_365_2822.n62 0.451587
R977 a_365_2822.n6 a_365_2822.n40 0.408833
R978 a_365_2822.n79 a_365_2822.n77 0.405391
R979 a_365_2822.n81 a_365_2822.n80 0.405391
R980 a_365_2822.n11 a_365_2822.n49 0.395292
R981 a_365_2822.n10 a_365_2822.n56 0.395292
R982 a_365_2822.n49 a_365_2822.n48 0.143208
R983 a_365_2822.n56 a_365_2822.n55 0.143208
R984 vcc.n30 vcc.n28 3045.88
R985 vcc.n32 vcc.n28 3045.88
R986 vcc.n32 vcc.n27 3045.88
R987 vcc.n30 vcc.n27 3045.88
R988 vcc.n77 vcc.n62 2704.62
R989 vcc.n77 vcc.n61 2699.48
R990 vcc.n74 vcc.n64 2372.5
R991 vcc.n74 vcc.n62 2327.31
R992 vcc.n56 vcc.n6 2089.41
R993 vcc.n53 vcc.n7 2089.41
R994 vcc.n45 vcc.n11 2089.41
R995 vcc.n48 vcc.n10 2089.41
R996 vcc.n41 vcc.n40 2089.41
R997 vcc.n38 vcc.n23 2089.41
R998 vcc.n76 vcc.t4 654.997
R999 vcc.t16 vcc.n62 616.96
R1000 vcc.n68 vcc.n67 599.49
R1001 vcc.t0 vcc.n27 538
R1002 vcc.n35 vcc.n24 524.801
R1003 vcc.t8 vcc.n28 524.534
R1004 vcc.n75 vcc.t16 519.274
R1005 vcc.n31 vcc.t8 441.339
R1006 vcc.n31 vcc.t0 427.875
R1007 vcc.n54 vcc.n6 426.346
R1008 vcc.n55 vcc.n7 426.346
R1009 vcc.n46 vcc.n45 426.346
R1010 vcc.n48 vcc.n47 426.346
R1011 vcc.n41 vcc.n21 426.346
R1012 vcc.n39 vcc.n38 426.346
R1013 vcc.t12 vcc.t4 387.817
R1014 vcc.n72 vcc.n71 298.611
R1015 vcc.n63 vcc.n61 268.716
R1016 vcc.n73 vcc.n66 253.067
R1017 vcc.n73 vcc.n72 248.246
R1018 vcc.n16 vcc.t15 231.286
R1019 vcc.n17 vcc.t11 231.286
R1020 vcc.n0 vcc.t7 231.286
R1021 vcc.n15 vcc.t9 231.273
R1022 vcc.n13 vcc.t1 231.272
R1023 vcc.n83 vcc.n1 202.453
R1024 vcc.n76 vcc.t2 196.603
R1025 vcc.t2 vcc.n75 168.089
R1026 vcc.n29 vcc.n26 128.857
R1027 vcc.n66 vcc.n65 118.645
R1028 vcc.n29 vcc.n24 103.353
R1029 vcc.n52 vcc.n4 101.719
R1030 vcc.n52 vcc.n51 82.4041
R1031 vcc.n43 vcc.n8 73.7015
R1032 vcc.n50 vcc.n8 72.4513
R1033 vcc.n65 vcc.n59 68.2096
R1034 vcc.n42 vcc.n12 64.5106
R1035 vcc.n36 vcc.n12 63.9989
R1036 vcc.n72 vcc.n62 61.6672
R1037 vcc.n67 vcc.t3 57.1305
R1038 vcc.n67 vcc.t17 57.1305
R1039 vcc.n66 vcc.n64 46.2505
R1040 vcc.n34 vcc.n33 44.5705
R1041 vcc.n33 vcc.n26 44.4238
R1042 vcc.n34 vcc.n25 40.7138
R1043 vcc.n25 vcc.n24 35.1619
R1044 vcc.n64 vcc.n63 33.6773
R1045 vcc.n27 vcc.n26 30.8799
R1046 vcc.n28 vcc.n25 30.8338
R1047 vcc.n38 vcc.n37 30.8338
R1048 vcc.n42 vcc.n41 30.8338
R1049 vcc.n45 vcc.n44 30.8338
R1050 vcc.n49 vcc.n48 30.8338
R1051 vcc.n6 vcc.n5 30.8338
R1052 vcc.n7 vcc.n4 30.8338
R1053 vcc.n65 vcc.n61 30.8338
R1054 vcc.n63 vcc.t12 29.2123
R1055 vcc.n1 vcc.t13 28.5655
R1056 vcc.n1 vcc.t5 28.5655
R1057 vcc.n58 vcc.n4 25.6005
R1058 vcc.n57 vcc.n56 23.1255
R1059 vcc.n11 vcc.n9 23.1255
R1060 vcc.n23 vcc.n12 23.1255
R1061 vcc.n40 vcc.n22 23.1255
R1062 vcc.n10 vcc.n8 23.1255
R1063 vcc.n53 vcc.n52 23.1255
R1064 vcc.n56 vcc.n55 18.2059
R1065 vcc.n47 vcc.n11 18.2059
R1066 vcc.n23 vcc.n21 18.2059
R1067 vcc.n40 vcc.n39 18.2059
R1068 vcc.n46 vcc.n10 18.2059
R1069 vcc.n54 vcc.n53 18.2059
R1070 vcc.n80 vcc.n59 14.5012
R1071 vcc.n79 vcc.n78 11.7493
R1072 vcc.n74 vcc.n73 11.563
R1073 vcc.n75 vcc.n74 11.563
R1074 vcc.n30 vcc.n29 10.8829
R1075 vcc.n31 vcc.n30 10.8829
R1076 vcc.n33 vcc.n32 10.8829
R1077 vcc.n32 vcc.n31 10.8829
R1078 vcc.n58 vcc.n57 9.4531
R1079 vcc.n51 vcc.n50 9.44208
R1080 vcc.n59 vcc.n58 9.35342
R1081 vcc.n79 vcc.n3 9.3005
R1082 vcc.n81 vcc.n80 9.3005
R1083 vcc.n44 vcc.n9 9.2534
R1084 vcc.n68 vcc 9.23317
R1085 vcc.n43 vcc.n42 9.22587
R1086 vcc.n57 vcc.n5 9.15071
R1087 vcc.n49 vcc.n9 9.1265
R1088 vcc.n37 vcc.n22 9.05594
R1089 vcc.n22 vcc.n20 8.90387
R1090 vcc.n36 vcc.n35 8.69513
R1091 vcc.n78 vcc.n77 7.4005
R1092 vcc.n77 vcc.n76 7.4005
R1093 vcc.t6 vcc.n54 4.71965
R1094 vcc.n55 vcc.t6 4.71965
R1095 vcc.t10 vcc.n46 4.71965
R1096 vcc.n47 vcc.t10 4.71965
R1097 vcc.n39 vcc.t14 4.71965
R1098 vcc.t14 vcc.n21 4.71965
R1099 vcc.n19 vcc.n14 3.76292
R1100 vcc.n82 vcc.n81 2.2505
R1101 vcc.n80 vcc.n79 1.2065
R1102 vcc.n78 vcc.n60 0.599649
R1103 vcc.n17 vcc.n0 0.53444
R1104 vcc.n16 vcc.n15 0.532497
R1105 vcc.n18 vcc.n17 0.492636
R1106 vcc.n70 vcc.n3 0.385704
R1107 vcc vcc.n83 0.331562
R1108 vcc.n13 vcc 0.293519
R1109 vcc.n71 vcc.n70 0.286982
R1110 vcc.n60 vcc.n2 0.239152
R1111 vcc.n44 vcc.n43 0.203427
R1112 vcc.n15 vcc.n14 0.177448
R1113 vcc.n82 vcc.n2 0.149902
R1114 vcc.n42 vcc.n20 0.109768
R1115 vcc.n69 vcc.n68 0.102498
R1116 vcc.n50 vcc.n49 0.0797079
R1117 vcc.n37 vcc.n36 0.0785488
R1118 vcc.n70 vcc.n69 0.0730806
R1119 vcc.n20 vcc.n19 0.0728582
R1120 vcc.n71 vcc.n60 0.064195
R1121 vcc.n14 vcc.n13 0.0593474
R1122 vcc.n51 vcc.n5 0.0480248
R1123 vcc.n18 vcc.n16 0.0423046
R1124 vcc.n81 vcc.n3 0.037915
R1125 vcc vcc.n0 0.0303013
R1126 vcc.n19 vcc.n18 0.0293462
R1127 vcc.n83 vcc.n82 0.0279096
R1128 vcc.n35 vcc.n34 0.0161098
R1129 vcc.n69 vcc.n2 0.000802663
R1130 vref.n4 vref.t0 231.292
R1131 vref.n3 vref.t4 85.987
R1132 vref.n2 vref.n0 71.7516
R1133 vref.n2 vref.n1 70.9453
R1134 vref.n0 vref.t3 17.4005
R1135 vref.n0 vref.t5 17.4005
R1136 vref.n1 vref.t1 17.4005
R1137 vref.n1 vref.t2 17.4005
R1138 vref.n4 vref.n3 1.0324
R1139 vref.n3 vref.n2 0.896828
R1140 vref vref.n4 0.408663
C0 a_4831_1286# a_3541_1286# 0.154516f
C1 a_3541_1286# BGR_BJT_stage1_0.vref0 0.011455f
C2 a_3541_1286# a_5031_1374# 1.04e-19
C3 vcc BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.50967f
C4 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2251_1286# 0.027078f
C5 vref vcc 0.285824f
C6 a_6121_1286# a_4831_1286# 0.154422f
C7 a_4831_1286# BGR_BJT_stage1_0.vref0 0.011274f
C8 a_3741_1374# vcc 0.034493f
C9 a_4831_1286# a_5031_1374# 1.53005f
C10 a_6121_1286# a_5031_1374# 0.10061f
C11 a_5031_1374# BGR_BJT_stage1_0.vref0 0.001349f
C12 vcc a_2451_1374# 0.034289f
C13 a_3741_1374# a_2251_1286# 1.04e-19
C14 a_2451_1374# a_2251_1286# 1.53765f
C15 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_3541_1286# 0.008224f
C16 a_3741_1374# a_3541_1286# 1.53781f
C17 a_3541_1286# a_2451_1374# 0.097608f
C18 a_4831_1286# BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.006534f
C19 a_6121_1286# BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.001655f
C20 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter BGR_BJT_stage1_0.vref0 16.430302f
C21 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_5031_1374# 1.25e-19
C22 vref a_4831_1286# 3.04e-19
C23 a_6121_1286# vref 1.65112f
C24 vref a_5031_1374# 0.036384f
C25 a_3741_1374# a_4831_1286# 0.098772f
C26 a_3741_1374# BGR_BJT_stage1_0.vref0 0.001621f
C27 a_3741_1374# a_5031_1374# 0.036353f
C28 a_2451_1374# BGR_BJT_stage1_0.vref0 0.03914f
C29 vcc a_2251_1286# 0.325293f
C30 vcc a_3541_1286# 0.319107f
C31 a_3541_1286# a_2251_1286# 0.154705f
C32 a_3741_1374# BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 1.25e-19
C33 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2451_1374# 0.002923f
C34 a_4831_1286# vcc 0.335825f
C35 a_6121_1286# vcc 0.368166f
C36 vcc BGR_BJT_stage1_0.vref0 0.05606f
C37 vcc a_5031_1374# 0.034455f
C38 a_3741_1374# a_2451_1374# 0.036353f
C39 a_2251_1286# BGR_BJT_stage1_0.vref0 0.114416f
C40 vref vss 0.942762f
C41 vcc vss 21.092445f
C42 a_5031_1374# vss 0.471213f
C43 a_3741_1374# vss 0.471213f
C44 a_2451_1374# vss 0.471599f
C45 a_6121_1286# vss 3.74418f
C46 a_4831_1286# vss 3.70955f
C47 a_3541_1286# vss 3.71022f
C48 a_2251_1286# vss 3.83691f
C49 BGR_BJT_stage1_0.vref0 vss 9.210018f
C50 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter vss 25.227676f
C51 vcc.t7 vss 0.009302f
C52 vcc.n0 vss 0.204711f
C53 vcc.t13 vss 0.002481f
C54 vcc.t5 vss 0.002481f
C55 vcc.n1 vss 0.005293f
C56 vcc.n2 vss 0.279031f
C57 vcc.n3 vss 0.031254f
C58 vcc.n4 vss 0.025624f
C59 vcc.n5 vss 0.08155f
C60 vcc.n6 vss 0.133363f
C61 vcc.n7 vss 0.133363f
C62 vcc.n8 vss 0.03008f
C63 vcc.n9 vss 0.129732f
C64 vcc.n10 vss 0.017637f
C65 vcc.n11 vss 0.017637f
C66 vcc.n12 vss 0.032126f
C67 vcc.t1 vss 0.0093f
C68 vcc.n13 vss 0.14272f
C69 vcc.n14 vss 0.159566f
C70 vcc.t15 vss 0.009302f
C71 vcc.t9 vss 0.009301f
C72 vcc.n15 vss 0.254353f
C73 vcc.n16 vss 0.208076f
C74 vcc.t11 vss 0.009302f
C75 vcc.n17 vss 0.349019f
C76 vcc.n18 vss 0.166659f
C77 vcc.n19 vss 0.544024f
C78 vcc.n20 vss 0.105461f
C79 vcc.n22 vss 0.12735f
C80 vcc.n23 vss 0.017637f
C81 vcc.n24 vss 0.032802f
C82 vcc.n25 vss 0.017469f
C83 vcc.n26 vss 0.10975f
C84 vcc.n27 vss 0.144915f
C85 vcc.n28 vss 0.140877f
C86 vcc.t0 vss 0.177019f
C87 vcc.t8 vss 0.176965f
C88 vcc.n29 vss 0.05086f
C89 vcc.n30 vss 0.025377f
C90 vcc.n31 vss 0.157827f
C91 vcc.n32 vss 0.025377f
C92 vcc.n33 vss 0.421347f
C93 vcc.n34 vss 0.068271f
C94 vcc.n35 vss 0.195811f
C95 vcc.n36 vss 0.216749f
C96 vcc.n37 vss 0.085226f
C97 vcc.n38 vss 0.133363f
C98 vcc.t14 vss 0.201185f
C99 vcc.n40 vss 0.017637f
C100 vcc.n41 vss 0.133363f
C101 vcc.n42 vss 0.228434f
C102 vcc.n43 vss 0.228718f
C103 vcc.n44 vss 0.082165f
C104 vcc.n45 vss 0.133363f
C105 vcc.t10 vss 0.201185f
C106 vcc.n48 vss 0.133363f
C107 vcc.n49 vss 0.082948f
C108 vcc.n50 vss 0.225245f
C109 vcc.n51 vss 0.223376f
C110 vcc.n52 vss 0.031431f
C111 vcc.n53 vss 0.017637f
C112 vcc.t6 vss 0.201185f
C113 vcc.n56 vss 0.017637f
C114 vcc.n57 vss 0.131204f
C115 vcc.n58 vss 0.164235f
C116 vcc.n59 vss 0.19526f
C117 vcc.n60 vss 0.09308f
C118 vcc.n61 vss 0.121712f
C119 vcc.n62 vss 0.165899f
C120 vcc.t4 vss 0.187615f
C121 vcc.t16 vss 0.206934f
C122 vcc.t12 vss 0.100507f
C123 vcc.n63 vss 0.044407f
C124 vcc.n64 vss 0.02929f
C125 vcc.n65 vss 0.020163f
C126 vcc.n66 vss 0.02929f
C127 vcc.t3 vss 0.001241f
C128 vcc.t17 vss 0.001241f
C129 vcc.n67 vss 0.002599f
C130 vcc.n68 vss 0.308488f
C131 vcc.n69 vss 0.059716f
C132 vcc.n70 vss 0.151717f
C133 vcc.n71 vss 0.394767f
C134 vcc.n72 vss 0.048834f
C135 vcc.n73 vss 0.039101f
C136 vcc.n74 vss 0.039101f
C137 vcc.n75 vss 0.124023f
C138 vcc.t2 vss 0.065802f
C139 vcc.n76 vss 0.153507f
C140 vcc.n77 vss 0.052409f
C141 vcc.n78 vss 0.090876f
C142 vcc.n79 vss 0.094691f
C143 vcc.n80 vss 0.11471f
C144 vcc.n81 vss 0.066281f
C145 vcc.n82 vss 0.104214f
C146 vcc.n83 vss 0.19103f
C147 a_365_2822.n0 vss 0.295573f
C148 a_365_2822.n1 vss 0.296251f
C149 a_365_2822.n2 vss 0.296328f
C150 a_365_2822.n3 vss 0.2939f
C151 a_365_2822.n4 vss 0.751854f
C152 a_365_2822.n5 vss 0.582261f
C153 a_365_2822.n6 vss 0.295548f
C154 a_365_2822.n7 vss 0.293282f
C155 a_365_2822.n8 vss 0.293737f
C156 a_365_2822.n9 vss 0.293309f
C157 a_365_2822.n10 vss 0.292124f
C158 a_365_2822.n11 vss 0.291156f
C159 a_365_2822.n12 vss 0.159721f
C160 a_365_2822.n13 vss 0.115661f
C161 a_365_2822.n14 vss 0.180826f
C162 a_365_2822.n15 vss 0.231328f
C163 a_365_2822.t47 vss 0.036484f
C164 a_365_2822.t30 vss 0.426788f
C165 a_365_2822.n16 vss 0.499268f
C166 a_365_2822.n17 vss 0.233812f
C167 a_365_2822.n18 vss 0.187249f
C168 a_365_2822.t8 vss 0.426145f
C169 a_365_2822.n19 vss 0.190828f
C170 a_365_2822.t36 vss 0.036484f
C171 a_365_2822.t19 vss 0.036484f
C172 a_365_2822.n20 vss 0.077885f
C173 a_365_2822.n21 vss 0.190696f
C174 a_365_2822.n22 vss 0.125951f
C175 a_365_2822.n23 vss 0.190841f
C176 a_365_2822.t18 vss 0.426145f
C177 a_365_2822.n24 vss 0.250942f
C178 a_365_2822.t26 vss 0.426145f
C179 a_365_2822.n25 vss 0.187651f
C180 a_365_2822.n26 vss 0.125933f
C181 a_365_2822.t27 vss 0.036484f
C182 a_365_2822.t45 vss 0.036484f
C183 a_365_2822.n27 vss 0.077885f
C184 a_365_2822.t32 vss 0.036484f
C185 a_365_2822.t9 vss 0.036484f
C186 a_365_2822.n28 vss 0.077885f
C187 a_365_2822.n29 vss 0.191394f
C188 a_365_2822.n30 vss 0.133088f
C189 a_365_2822.n31 vss 0.195738f
C190 a_365_2822.t10 vss 0.426145f
C191 a_365_2822.n32 vss 0.191935f
C192 a_365_2822.t0 vss 0.426145f
C193 a_365_2822.n33 vss 0.189447f
C194 a_365_2822.t28 vss 0.426145f
C195 a_365_2822.n34 vss 0.19169f
C196 a_365_2822.t11 vss 0.036484f
C197 a_365_2822.t33 vss 0.036484f
C198 a_365_2822.n35 vss 0.077885f
C199 a_365_2822.t40 vss 0.036484f
C200 a_365_2822.t29 vss 0.036484f
C201 a_365_2822.n36 vss 0.077885f
C202 a_365_2822.t17 vss 0.036484f
C203 a_365_2822.t42 vss 0.036484f
C204 a_365_2822.n37 vss 0.078094f
C205 a_365_2822.t16 vss 0.426145f
C206 a_365_2822.n38 vss 0.193366f
C207 a_365_2822.n39 vss 0.127361f
C208 a_365_2822.n40 vss 0.109271f
C209 a_365_2822.n41 vss 0.125951f
C210 a_365_2822.n42 vss 0.250961f
C211 a_365_2822.n43 vss 0.283641f
C212 a_365_2822.n44 vss 0.184132f
C213 a_365_2822.n45 vss 0.125976f
C214 a_365_2822.t25 vss 0.036484f
C215 a_365_2822.t43 vss 0.036484f
C216 a_365_2822.n46 vss 0.077937f
C217 a_365_2822.t39 vss 0.036484f
C218 a_365_2822.t3 vss 0.036484f
C219 a_365_2822.n47 vss 0.077939f
C220 a_365_2822.n48 vss 0.223243f
C221 a_365_2822.n49 vss 0.074968f
C222 a_365_2822.t2 vss 0.426145f
C223 a_365_2822.n50 vss 0.187249f
C224 a_365_2822.t14 vss 0.426145f
C225 a_365_2822.n51 vss 0.190252f
C226 a_365_2822.n52 vss 0.115915f
C227 a_365_2822.t15 vss 0.036484f
C228 a_365_2822.t44 vss 0.036484f
C229 a_365_2822.n53 vss 0.077937f
C230 a_365_2822.t41 vss 0.036484f
C231 a_365_2822.t7 vss 0.036484f
C232 a_365_2822.n54 vss 0.077937f
C233 a_365_2822.n55 vss 0.223409f
C234 a_365_2822.n56 vss 0.073836f
C235 a_365_2822.t12 vss 0.426781f
C236 a_365_2822.n57 vss 0.509608f
C237 a_365_2822.t37 vss 0.036484f
C238 a_365_2822.t13 vss 0.036484f
C239 a_365_2822.n58 vss 0.077937f
C240 a_365_2822.n59 vss 0.279619f
C241 a_365_2822.t5 vss 0.036484f
C242 a_365_2822.t35 vss 0.036484f
C243 a_365_2822.n60 vss 0.077937f
C244 a_365_2822.n61 vss 0.125933f
C245 a_365_2822.t4 vss 0.426145f
C246 a_365_2822.n62 vss 0.194649f
C247 a_365_2822.n63 vss 0.19363f
C248 a_365_2822.t6 vss 0.426145f
C249 a_365_2822.n64 vss 0.23377f
C250 a_365_2822.n65 vss 0.159699f
C251 a_365_2822.n66 vss 0.173683f
C252 a_365_2822.n67 vss 0.250389f
C253 a_365_2822.n68 vss 0.125951f
C254 a_365_2822.t34 vss 0.036484f
C255 a_365_2822.t1 vss 0.036484f
C256 a_365_2822.n69 vss 0.077885f
C257 a_365_2822.t21 vss 0.036484f
C258 a_365_2822.t46 vss 0.036484f
C259 a_365_2822.n70 vss 0.077885f
C260 a_365_2822.t20 vss 0.426145f
C261 a_365_2822.n71 vss 0.191677f
C262 a_365_2822.n72 vss 0.125933f
C263 a_365_2822.n73 vss 0.125952f
C264 a_365_2822.n74 vss 0.250976f
C265 a_365_2822.n75 vss 0.173683f
C266 a_365_2822.n76 vss 0.159699f
C267 a_365_2822.n77 vss 0.243651f
C268 a_365_2822.n78 vss 0.151692f
C269 a_365_2822.n79 vss 0.197087f
C270 a_365_2822.t24 vss 0.426145f
C271 a_365_2822.n80 vss 0.208755f
C272 a_365_2822.t22 vss 0.426145f
C273 a_365_2822.n81 vss 0.209523f
C274 a_365_2822.n82 vss 0.151723f
C275 a_365_2822.t38 vss 0.036484f
C276 a_365_2822.t23 vss 0.036484f
C277 a_365_2822.n83 vss 0.077937f
C278 a_365_2822.n84 vss 0.077937f
C279 a_365_2822.t31 vss 0.036484f
C280 BGR_BJT_stage1_0.vref0.n0 vss 1.13777f
C281 BGR_BJT_stage1_0.vref0.t6 vss 0.079462f
C282 BGR_BJT_stage1_0.vref0.t2 vss 0.079462f
C283 BGR_BJT_stage1_0.vref0.n1 vss 0.255115f
C284 BGR_BJT_stage1_0.vref0.t1 vss 0.079462f
C285 BGR_BJT_stage1_0.vref0.t19 vss 0.079462f
C286 BGR_BJT_stage1_0.vref0.n2 vss 0.255115f
C287 BGR_BJT_stage1_0.vref0.t11 vss 0.079462f
C288 BGR_BJT_stage1_0.vref0.t25 vss 0.079462f
C289 BGR_BJT_stage1_0.vref0.n3 vss 0.255115f
C290 BGR_BJT_stage1_0.vref0.t14 vss 0.079462f
C291 BGR_BJT_stage1_0.vref0.t3 vss 0.079462f
C292 BGR_BJT_stage1_0.vref0.n4 vss 0.255115f
C293 BGR_BJT_stage1_0.vref0.t27 vss 0.079462f
C294 BGR_BJT_stage1_0.vref0.t10 vss 0.079462f
C295 BGR_BJT_stage1_0.vref0.n5 vss 0.265118f
C296 BGR_BJT_stage1_0.vref0.n6 vss 1.61061f
C297 BGR_BJT_stage1_0.vref0.t22 vss 0.079462f
C298 BGR_BJT_stage1_0.vref0.t21 vss 0.079462f
C299 BGR_BJT_stage1_0.vref0.n7 vss 0.255115f
C300 BGR_BJT_stage1_0.vref0.n8 vss 0.934734f
C301 BGR_BJT_stage1_0.vref0.n9 vss 0.934734f
C302 BGR_BJT_stage1_0.vref0.n10 vss 0.934734f
C303 BGR_BJT_stage1_0.vref0.n11 vss 0.91495f
C304 BGR_BJT_stage1_0.vref0.t30 vss 0.079462f
C305 BGR_BJT_stage1_0.vref0.t13 vss 0.079462f
C306 BGR_BJT_stage1_0.vref0.n12 vss 0.255115f
C307 BGR_BJT_stage1_0.vref0.t9 vss 0.079462f
C308 BGR_BJT_stage1_0.vref0.t32 vss 0.079462f
C309 BGR_BJT_stage1_0.vref0.n13 vss 0.254999f
C310 BGR_BJT_stage1_0.vref0.t12 vss 0.079462f
C311 BGR_BJT_stage1_0.vref0.t4 vss 0.079462f
C312 BGR_BJT_stage1_0.vref0.n14 vss 0.278374f
C313 BGR_BJT_stage1_0.vref0.t28 vss 0.079462f
C314 BGR_BJT_stage1_0.vref0.t7 vss 0.079462f
C315 BGR_BJT_stage1_0.vref0.n15 vss 0.254679f
C316 BGR_BJT_stage1_0.vref0.n16 vss 1.71688f
C317 BGR_BJT_stage1_0.vref0.t8 vss 0.079462f
C318 BGR_BJT_stage1_0.vref0.t24 vss 0.079462f
C319 BGR_BJT_stage1_0.vref0.n17 vss 0.254679f
C320 BGR_BJT_stage1_0.vref0.n18 vss 0.925607f
C321 BGR_BJT_stage1_0.vref0.t29 vss 0.079462f
C322 BGR_BJT_stage1_0.vref0.t15 vss 0.079462f
C323 BGR_BJT_stage1_0.vref0.n19 vss 0.254679f
C324 BGR_BJT_stage1_0.vref0.n20 vss 0.925607f
C325 BGR_BJT_stage1_0.vref0.t20 vss 0.079462f
C326 BGR_BJT_stage1_0.vref0.t5 vss 0.079462f
C327 BGR_BJT_stage1_0.vref0.n21 vss 0.254679f
C328 BGR_BJT_stage1_0.vref0.n22 vss 0.925607f
C329 BGR_BJT_stage1_0.vref0.t31 vss 0.079462f
C330 BGR_BJT_stage1_0.vref0.t17 vss 0.079462f
C331 BGR_BJT_stage1_0.vref0.n23 vss 0.254679f
C332 BGR_BJT_stage1_0.vref0.n24 vss 0.925607f
C333 BGR_BJT_stage1_0.vref0.t16 vss 0.079462f
C334 BGR_BJT_stage1_0.vref0.t23 vss 0.079462f
C335 BGR_BJT_stage1_0.vref0.n25 vss 0.254679f
C336 BGR_BJT_stage1_0.vref0.n26 vss 0.925607f
C337 BGR_BJT_stage1_0.vref0.t26 vss 0.079462f
C338 BGR_BJT_stage1_0.vref0.t18 vss 0.079462f
C339 BGR_BJT_stage1_0.vref0.n27 vss 0.254679f
C340 BGR_BJT_stage1_0.vref0.n28 vss 1.44007f
C341 BGR_BJT_stage1_0.vref0.n29 vss 1.30818f
C342 BGR_BJT_stage1_0.vref0.t0 vss 0.077176f
C343 BGR_BJT_stage1_0.vr.n0 vss 3.30312f
C344 BGR_BJT_stage1_0.vr.n1 vss 6.26335f
C345 BGR_BJT_stage1_0.vr.n2 vss 3.66726f
C346 BGR_BJT_stage2_0.vr vss 1.01868f
C347 BGR_BJT_stage1_0.vr.t26 vss 0.607494f
C348 BGR_BJT_stage1_0.vr.t24 vss 0.584182f
C349 BGR_BJT_stage1_0.vr.n3 vss 1.65172f
C350 BGR_BJT_stage1_0.vr.t21 vss 0.584182f
C351 BGR_BJT_stage1_0.vr.n4 vss 0.975793f
C352 BGR_BJT_stage1_0.vr.t23 vss 0.584182f
C353 BGR_BJT_stage1_0.vr.n5 vss 0.974491f
C354 BGR_BJT_stage1_0.vr.t20 vss 0.584182f
C355 BGR_BJT_stage1_0.vr.t25 vss 0.303271f
C356 BGR_BJT_stage1_0.vr.t1 vss 0.025822f
C357 BGR_BJT_stage1_0.vr.t3 vss 0.025857f
C358 BGR_BJT_stage1_0.vr.t2 vss 0.45849f
C359 BGR_BJT_stage1_0.vr.t8 vss 0.275911f
C360 BGR_BJT_stage1_0.vr.t18 vss 0.054718f
C361 BGR_BJT_stage1_0.vr.t11 vss 0.054718f
C362 BGR_BJT_stage1_0.vr.n6 vss 0.207857f
C363 BGR_BJT_stage1_0.vr.t6 vss 0.054718f
C364 BGR_BJT_stage1_0.vr.t14 vss 0.054718f
C365 BGR_BJT_stage1_0.vr.n7 vss 0.207857f
C366 BGR_BJT_stage1_0.vr.t15 vss 0.054718f
C367 BGR_BJT_stage1_0.vr.t12 vss 0.054718f
C368 BGR_BJT_stage1_0.vr.n8 vss 0.207857f
C369 BGR_BJT_stage1_0.vr.t19 vss 0.301217f
C370 BGR_BJT_stage1_0.vr.t13 vss 0.054718f
C371 BGR_BJT_stage1_0.vr.t10 vss 0.054718f
C372 BGR_BJT_stage1_0.vr.n9 vss 0.207857f
C373 BGR_BJT_stage1_0.vr.t16 vss 0.054718f
C374 BGR_BJT_stage1_0.vr.t7 vss 0.054718f
C375 BGR_BJT_stage1_0.vr.n10 vss 0.207857f
C376 BGR_BJT_stage1_0.vr.t9 vss 0.054718f
C377 BGR_BJT_stage1_0.vr.t5 vss 0.054718f
C378 BGR_BJT_stage1_0.vr.n11 vss 0.207857f
C379 BGR_BJT_stage1_0.vr.t4 vss 0.054718f
C380 BGR_BJT_stage1_0.vr.t17 vss 0.054718f
C381 BGR_BJT_stage1_0.vr.n12 vss 0.236074f
C382 BGR_BJT_stage1_0.vr.t0 vss 0.45849f
C383 BGR_BJT_stage1_0.vr.t22 vss 0.30303f
C384 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 vss 0.072341f
C385 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 vss 0.122613f
C386 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 vss 0.215544f
C387 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 vss 0.480953f
C388 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 vss 0.479714f
C389 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 vss 1.17298f
C390 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 vss 0.305899f
C391 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 vss 0.47876f
C392 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 vss 0.234546f
C393 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 vss 0.471294f
C394 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 vss 0.47876f
C395 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 vss 0.471294f
C396 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 vss 0.47876f
C397 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 vss 0.470848f
C398 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 vss 0.47876f
C399 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 vss 0.119506f
C400 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 vss 0.391762f
C401 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 vss 0.208072f
C402 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 vss 0.305783f
C403 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 vss 0.479542f
C404 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 vss 0.222367f
C405 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 vss 0.474879f
C406 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 vss 0.47876f
C407 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 vss 0.474879f
C408 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 vss 0.47876f
C409 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 vss 0.472824f
C410 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 vss 0.47876f
C411 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 vss 0.114778f
C412 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 vss 0.358618f
C413 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 vss 0.171563f
C414 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 vss 0.305632f
C415 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 vss 0.47876f
C416 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 vss 0.235085f
C417 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 vss 0.471837f
C418 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 vss 0.47876f
C419 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 vss 0.471837f
C420 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 vss 0.47876f
C421 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 vss 0.471737f
C422 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 vss 0.47876f
C423 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 vss 0.11683f
C424 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 vss 0.392517f
C425 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 vss 0.175671f
C426 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 vss 0.305654f
C427 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 vss 0.479614f
C428 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 vss 0.233152f
C429 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 vss 0.470751f
C430 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 vss 0.47876f
C431 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 vss 0.470751f
C432 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 vss 0.47876f
C433 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 vss 0.471056f
C434 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 vss 0.47876f
C435 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 vss 0.119137f
C436 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 vss 0.357782f
C437 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 vss 0.171642f
C438 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 vss 0.306196f
C439 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 vss 0.47876f
C440 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 vss 0.231876f
C441 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 vss 0.471573f
C442 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 vss 0.47876f
C443 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 vss 0.471573f
C444 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 vss 0.47876f
C445 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 vss 0.467455f
C446 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 vss 0.47876f
C447 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 vss 0.124281f
C448 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 vss 0.392522f
C449 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 vss 0.175671f
C450 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 vss 0.158535f
C451 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 vss 0.47876f
C452 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 vss 0.47876f
C453 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 vss 0.304891f
C454 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 vss 0.158873f
C455 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 vss 0.478766f
C456 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 vss 0.29558f
C457 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 vss 0.280101f
C458 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 vss 0.461265f
C459 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 vss 0.301638f
C460 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 vss 0.282184f
C461 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 vss 0.47876f
C462 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 vss 0.208844f
C463 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 vss 0.172117f
C464 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 vss 0.305976f
C465 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 vss 0.47876f
C466 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 vss 0.22879f
C467 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 vss 0.474578f
C468 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 vss 0.47876f
C469 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 vss 0.474578f
C470 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 vss 0.47876f
C471 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 vss 0.473804f
C472 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 vss 0.47876f
C473 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 vss 0.113869f
C474 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 vss 0.395959f
C475 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 vss 0.1767f
C476 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 vss 0.294557f
C477 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 vss 0.47876f
C478 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 vss 0.283413f
C479 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 vss 0.47876f
C480 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 vss 0.443727f
C481 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 vss 0.195453f
C482 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 vss 0.373404f
C483 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 vss 0.49099f
C484 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 vss 0.122613f
C485 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 vss 0.041314f
C486 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 vss 0.041318f
C487 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 vss 1.05832f
C488 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 vss 0.709094f
C489 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 vss 0.50264f
C490 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 vss 0.160856f
C491 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 vss 0.201533f
C492 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 vss 0.215544f
C493 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 vss 0.110351f
C494 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 vss 0.110351f
C495 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 vss 0.122613f
C496 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 vss 0.109327f
C497 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 vss 0.108125f
C498 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 vss 0.215049f
C499 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 vss 0.216251f
C500 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 vss 0.063674f
C501 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 vss 0.215593f
C502 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 vss 0.315796f
C503 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 vss 0.473909f
C504 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 vss 0.215544f
C505 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 vss 0.077246f
.ends

