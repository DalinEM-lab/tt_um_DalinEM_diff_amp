* NGSPICE file created from tt_um_DalinEM_diff_amp.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_L4HHUA a_n258_n100# a_n200_n197# a_200_n100# w_n294_n200#
X0 a_200_n100# a_n200_n197# a_n258_n100# w_n294_n200# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_LH3874 a_100_n100# a_n158_n100# a_n100_n188# VSUBS
X0 a_100_n100# a_n100_n188# a_n158_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_QCP9T2 a_n258_n100# a_n200_n197# a_200_n100# w_n294_n200#
X0 a_200_n100# a_n200_n197# a_n258_n100# w_n294_n200# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_Q4S9T2 a_n258_n100# w_n396_n319# a_n200_n197#
+ a_200_n100#
X0 a_200_n100# a_n200_n197# a_n258_n100# w_n396_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt BGR_BJT_stage2 vcc vss vref vref0 vr
XXM12 vcc vr vref vcc sky130_fd_pr__pfet_01v8_lvt_L4HHUA
XXM23 vref m1_4340_877# m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM13 m1_846_923# m1_971_877# m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM24 m1_4340_877# vref m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM15 m1_3032_877# m1_2136_923# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM16 m1_2136_923# m1_846_923# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM17 vcc vr m1_4340_877# vcc sky130_fd_pr__pfet_01v8_lvt_QCP9T2
XXM18 m1_4340_877# vref m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM19 vref m1_2136_923# m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM1 m1_n444_923# m1_75_833# m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM2 m1_75_833# m1_n444_923# m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM3 m1_n444_923# m1_75_833# m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM4 m1_n444_923# vref0 m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM5 m1_75_833# m1_n444_923# m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM6 m1_846_923# m1_n444_923# m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
Xsky130_fd_pr__nfet_01v8_lvt_LH3874_0 vref m1_4340_877# m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM7 m1_971_877# m1_846_923# m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM8 m1_846_923# m1_971_877# m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM9 m1_971_877# m1_846_923# m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
Xsky130_fd_pr__pfet_01v8_lvt_Q4S9T2_0 vcc vcc vr m1_3032_877# sky130_fd_pr__pfet_01v8_lvt_Q4S9T2
Xsky130_fd_pr__pfet_01v8_lvt_Q4S9T2_1 vcc vcc vr m1_75_833# sky130_fd_pr__pfet_01v8_lvt_Q4S9T2
XXM20 m1_2136_923# m1_3032_877# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM21 m1_3032_877# m1_2136_923# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM11 vcc vcc vr m1_971_877# sky130_fd_pr__pfet_01v8_lvt_Q4S9T2
XXM22 m1_2136_923# m1_3032_877# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2 a_100_n400# a_n158_n400# a_n100_n488# VSUBS
X0 a_100_n400# a_n100_n488# a_n158_n400# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_KLHH7J a_n200_n147# a_n258_n50# a_200_n50# w_n294_n150#
X0 a_200_n50# a_n200_n147# a_n258_n50# w_n294_n150# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_QCPJZY a_n100_n197# a_100_n100# w_n194_n200# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n194_n200# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
.ends

.subckt BGR_BJT_stage1 vcc vref0 vr vss
XXM12 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM23 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM34 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM45 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM14 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM24 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM25 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM35 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM36 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM46 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM47 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM15 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM26 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM37 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM48 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM16 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM27 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM38 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM49 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM17 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM28 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM39 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM18 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM29 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM19 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM1 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM2 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM3 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM4 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM5 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM6 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM7 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM8 vr vr vcc vcc sky130_fd_pr__pfet_01v8_lvt_KLHH7J
XXM9 vr vcc vcc sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter sky130_fd_pr__pfet_01v8_lvt_QCPJZY
Xsky130_fd_pr__nfet_01v8_lvt_UZ3GQ2_0 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__pfet_01v8_lvt_KLHH7J_0 vr vcc vr vcc sky130_fd_pr__pfet_01v8_lvt_KLHH7J
XXM50 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__pfet_01v8_lvt_QCPJZY_0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
+ vcc vcc sky130_fd_pr__pfet_01v8_lvt_QCPJZY
XXM40 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
+ vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXM30 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM41 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM20 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM31 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM42 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM10 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM21 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM32 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM43 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM11 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM22 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM33 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM44 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
.ends

.subckt BGR_BJT_vref vref vcc vss
XBGR_BJT_stage2_0 vcc vss vref BGR_BJT_stage2_0/vref0 BGR_BJT_stage2_0/vr BGR_BJT_stage2
XBGR_BJT_stage1_0 vcc BGR_BJT_stage2_0/vref0 BGR_BJT_stage2_0/vr vss BGR_BJT_stage1
.ends

.subckt OTA_vref_stage2 vcc vss vb vref0 vr vb1
XXM12 vcc vr vb vcc sky130_fd_pr__pfet_01v8_lvt_L4HHUA
XXM23 vb m1_4340_877# m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM13 vb1 m1_971_877# m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM24 m1_4340_877# vb m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM15 m1_3032_877# m1_2136_923# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM16 m1_2136_923# vb1 m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM17 vcc vr m1_4340_877# vcc sky130_fd_pr__pfet_01v8_lvt_QCP9T2
XXM18 m1_4340_877# vb m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM19 vb m1_2136_923# m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM1 m1_n444_923# m1_75_833# m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM2 m1_75_833# m1_n444_923# m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM3 m1_n444_923# m1_75_833# m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM4 m1_n444_923# vref0 m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM5 m1_75_833# m1_n444_923# m1_75_833# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM6 vb1 m1_n444_923# m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
Xsky130_fd_pr__nfet_01v8_lvt_LH3874_0 vb m1_4340_877# m1_4340_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM7 m1_971_877# vb1 m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM8 vb1 m1_971_877# m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM9 m1_971_877# vb1 m1_971_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
Xsky130_fd_pr__pfet_01v8_lvt_Q4S9T2_0 vcc vcc vr m1_3032_877# sky130_fd_pr__pfet_01v8_lvt_Q4S9T2
Xsky130_fd_pr__pfet_01v8_lvt_Q4S9T2_1 vcc vcc vr m1_75_833# sky130_fd_pr__pfet_01v8_lvt_Q4S9T2
XXM20 m1_2136_923# m1_3032_877# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM21 m1_3032_877# m1_2136_923# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
XXM11 vcc vcc vr m1_971_877# sky130_fd_pr__pfet_01v8_lvt_Q4S9T2
XXM22 m1_2136_923# m1_3032_877# m1_3032_877# vss sky130_fd_pr__nfet_01v8_lvt_LH3874
.ends

.subckt OTA_vref_stage1 vcc vref0 vr vss
XXM12 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM23 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM34 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM45 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM14 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM24 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM25 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM35 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM36 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM46 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM47 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM15 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM26 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM37 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM48 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM16 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM27 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM38 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM49 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM17 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM28 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM39 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM18 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM29 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM19 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM1 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM2 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM3 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM4 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM5 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM6 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM7 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM8 vr vr vcc vcc sky130_fd_pr__pfet_01v8_lvt_KLHH7J
XXM9 vr vcc vcc sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter sky130_fd_pr__pfet_01v8_lvt_QCPJZY
Xsky130_fd_pr__nfet_01v8_lvt_UZ3GQ2_0 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__pfet_01v8_lvt_KLHH7J_0 vr vcc vr vcc sky130_fd_pr__pfet_01v8_lvt_KLHH7J
XXM50 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__pfet_01v8_lvt_QCPJZY_0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
+ vcc vcc sky130_fd_pr__pfet_01v8_lvt_QCPJZY
XXM40 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
+ vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXM30 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM41 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM20 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM31 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM42 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM10 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM21 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM32 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM43 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM11 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM22 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM33 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM44 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
.ends

.subckt OTA_vref vb vb1 vcc vss
XOTA_vref_stage2_0 vcc vss vb OTA_vref_stage2_0/vref0 OTA_vref_stage2_0/vr vb1 OTA_vref_stage2
XOTA_vref_stage1_0 vcc OTA_vref_stage2_0/vref0 OTA_vref_stage2_0/vr vss OTA_vref_stage1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_NH7ZMU a_n190_n1597# a_190_n1500# w_n284_n1600#
+ a_n248_n1500#
X0 a_190_n1500# a_n190_n1597# a_n248_n1500# w_n284_n1600# sky130_fd_pr__pfet_01v8_lvt ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=1.9
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AR4WA2 a_n940_n238# a_940_n150# a_n998_n150# VSUBS
X0 a_940_n150# a_n940_n238# a_n998_n150# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=9.4
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_Q9T44L a_n35_n516# a_n165_n646# a_n35_84#
X0 a_n35_84# a_n35_n516# a_n165_n646# sky130_fd_pr__res_xhigh_po_0p35 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_6JHA76 a_n29_n700# w_n1003_n919# a_n865_n700# a_29_n797#
+ a_n807_n797# a_807_n700# a_n447_n700# a_n389_n797# a_389_n700# a_447_n797#
X0 a_807_n700# a_447_n797# a_389_n700# w_n1003_n919# sky130_fd_pr__pfet_01v8 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=1.8
X1 a_n447_n700# a_n807_n797# a_n865_n700# w_n1003_n919# sky130_fd_pr__pfet_01v8 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=1.8
X2 a_n29_n700# a_n389_n797# a_n447_n700# w_n1003_n919# sky130_fd_pr__pfet_01v8 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1.8
X3 a_389_n700# a_29_n797# a_n29_n700# w_n1003_n919# sky130_fd_pr__pfet_01v8 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1.8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_V6F9HY c1_n2146_n2000# m3_n2186_n2040#
X0 c1_n2146_n2000# m3_n2186_n2040# sky130_fd_pr__cap_mim_m3_1 l=20 w=20
.ends

.subckt OTA_stage2 vcc vss vo vd1 vd2 vb1
XXM12 vd1 vo vcc m1_7238_n2948# sky130_fd_pr__pfet_01v8_lvt_NH7ZMU
XXM15 m1_6804_n972# m1_6804_n972# vss vss sky130_fd_pr__nfet_01v8_lvt_AR4WA2
XXM16 m1_6804_n972# m1_6804_n972# vss vss sky130_fd_pr__nfet_01v8_lvt_AR4WA2
XXM17 m1_6804_n972# vss m1_6804_n972# vss sky130_fd_pr__nfet_01v8_lvt_AR4WA2
XXM18 m1_6804_n972# vss vo vss sky130_fd_pr__nfet_01v8_lvt_AR4WA2
XXM19 m1_6804_n972# vss vo vss sky130_fd_pr__nfet_01v8_lvt_AR4WA2
XXR34 vo vss m1_14583_n1665# sky130_fd_pr__res_xhigh_po_0p35_Q9T44L
XXM3 m1_7238_n2948# vcc m1_7238_n2948# vb1 vb1 m1_7238_n2948# vcc vb1 vcc vb1 sky130_fd_pr__pfet_01v8_6JHA76
XXM4 vd2 m1_6804_n972# vcc m1_7238_n2948# sky130_fd_pr__pfet_01v8_lvt_NH7ZMU
XXM5 vd2 m1_7238_n2948# vcc m1_6804_n972# sky130_fd_pr__pfet_01v8_lvt_NH7ZMU
XXM7 vd2 m1_7238_n2948# vcc m1_6804_n972# sky130_fd_pr__pfet_01v8_lvt_NH7ZMU
XXM8 vd1 m1_7238_n2948# vcc vo sky130_fd_pr__pfet_01v8_lvt_NH7ZMU
XXM9 m1_6804_n972# vss m1_6804_n972# vss sky130_fd_pr__nfet_01v8_lvt_AR4WA2
XXC1 m1_14583_n1665# vd1 sky130_fd_pr__cap_mim_m3_1_V6F9HY
Xsky130_fd_pr__pfet_01v8_lvt_NH7ZMU_0 vd1 m1_7238_n2948# vcc vo sky130_fd_pr__pfet_01v8_lvt_NH7ZMU
Xsky130_fd_pr__pfet_01v8_lvt_NH7ZMU_1 vd1 vo vcc m1_7238_n2948# sky130_fd_pr__pfet_01v8_lvt_NH7ZMU
Xsky130_fd_pr__nfet_01v8_lvt_AR4WA2_0 m1_6804_n972# vo vss vss sky130_fd_pr__nfet_01v8_lvt_AR4WA2
XXM10 m1_6804_n972# vo vss vss sky130_fd_pr__nfet_01v8_lvt_AR4WA2
XXM11 vd2 m1_6804_n972# vcc m1_7238_n2948# sky130_fd_pr__pfet_01v8_lvt_NH7ZMU
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_58FN7G a_n1800_n277# a_1800_n180# a_n1858_n180#
+ w_n1894_n280#
X0 a_1800_n180# a_n1800_n277# a_n1858_n180# w_n1894_n280# sky130_fd_pr__pfet_01v8_lvt ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=18
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_59CFV9 a_1200_n600# a_n1258_n600# a_n1200_n688#
+ VSUBS
X0 a_1200_n600# a_n1200_n688# a_n1258_n600# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=12
.ends

.subckt sky130_fd_pr__nfet_01v8_Q93DRV a_n558_n300# a_n500_n388# a_n660_n474# a_500_n300#
X0 a_500_n300# a_n500_n388# a_n558_n300# a_n660_n474# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=5
.ends

.subckt OTA_stage1 vd1 vin_p vin_n vb vcc vss vd2
Xsky130_fd_pr__pfet_01v8_lvt_58FN7G_0 vd2 vd1 vcc vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM1 m1_11317_n793# vd2 vin_p vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM2 m1_11317_n793# vd1 vin_n vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM3 vss vb vss m1_11317_n793# sky130_fd_pr__nfet_01v8_Q93DRV
XXM4 vd2 vcc vd1 vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM5 vd2 vcc vd2 vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM6 vd2 vd2 vcc vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
Xsky130_fd_pr__nfet_01v8_lvt_59CFV9_0 vd1 m1_11317_n793# vin_n vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM8 vd2 m1_11317_n793# vin_p vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
.ends

.subckt x2_OTA vo vin_p vin_n vss vcc
XOTA_vref_0 OTA_vref_0/vb OTA_vref_0/vb1 vcc vss OTA_vref
XOTA_stage2_0 vcc vss vo OTA_stage2_0/vd1 OTA_stage2_0/vd2 OTA_vref_0/vb1 OTA_stage2
XOTA_stage1_0 OTA_stage2_0/vd1 vin_p vin_n OTA_vref_0/vb vcc vss OTA_stage2_0/vd2
+ OTA_stage1
.ends

.subckt diff_final_v0 vout vin_p vin_n vb vcc vss
Xsky130_fd_pr__pfet_01v8_lvt_58FN7G_0 m1_15336_1751# vout vcc vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM1 m1_11317_n793# m1_15336_1751# vin_p vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM2 m1_11317_n793# vout vin_n vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM3 vss vb vss m1_11317_n793# sky130_fd_pr__nfet_01v8_Q93DRV
XXM4 m1_15336_1751# vcc vout vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM5 m1_15336_1751# vcc m1_15336_1751# vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
XXM6 m1_15336_1751# m1_15336_1751# vcc vcc sky130_fd_pr__pfet_01v8_lvt_58FN7G
Xsky130_fd_pr__nfet_01v8_lvt_59CFV9_0 vout m1_11317_n793# vin_n vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
XXM8 m1_15336_1751# m1_11317_n793# vin_p vss sky130_fd_pr__nfet_01v8_lvt_59CFV9
.ends

.subckt tt_um_DalinEM_diff_amp clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] VDPWR VGND
XBGR_BJT_vref_0 ua[5] VDPWR VGND BGR_BJT_vref
X2_OTA_0 ua[0] ua[2] ua[3] VGND VDPWR x2_OTA
Xdiff_final_v0_0 ua[1] ua[2] ua[3] ua[4] VDPWR VGND diff_final_v0
.ends

