magic
tech sky130A
magscale 1 2
timestamp 1738634814
<< nwell >>
rect 5611 -2535 7764 -1863
rect 6853 -2537 7764 -2535
<< pwell >>
rect 5516 949 12358 2193
rect 5516 945 7676 949
rect 7708 945 12358 949
rect 5516 899 12358 945
rect 5516 896 7674 899
rect 7707 896 12358 899
rect 5516 -921 12358 896
<< psubdiff >>
rect 5630 2019 5690 2053
rect 12146 2019 12206 2053
rect 5630 1993 5664 2019
rect 5630 -742 5664 -716
rect 12172 1993 12206 2019
rect 12172 -742 12206 -716
rect 5630 -776 5690 -742
rect 12146 -776 12206 -742
<< nsubdiff >>
rect 5740 -1940 5800 -1906
rect 6838 -1940 6898 -1906
rect 5740 -1966 5774 -1940
rect 5740 -2350 5774 -2324
rect 6864 -1966 6898 -1940
rect 6864 -2350 6898 -2324
rect 5740 -2384 5800 -2350
rect 6838 -2384 6898 -2350
<< psubdiffcont >>
rect 5690 2019 12146 2053
rect 5630 -716 5664 1993
rect 12172 -716 12206 1993
rect 5690 -776 12146 -742
<< nsubdiffcont >>
rect 5800 -1940 6838 -1906
rect 5740 -2324 5774 -1966
rect 6864 -2324 6898 -1966
rect 5800 -2384 6838 -2350
<< locali >>
rect 5511 2190 12229 2268
rect 5511 2016 5614 2190
rect 12192 2016 12229 2190
rect 5511 1993 12229 2016
rect 5511 1907 5630 1993
rect 5598 -716 5630 1907
rect 5664 1907 12172 1993
rect 5664 -706 5690 1907
rect 12113 -699 12172 1907
rect 5850 -706 12172 -699
rect 5664 -716 12172 -706
rect 12206 -716 12229 1993
rect 5598 -742 12229 -716
rect 5598 -776 5690 -742
rect 12146 -751 12229 -742
rect 5598 -863 5807 -776
rect 12148 -863 12229 -751
rect 5598 -907 12229 -863
rect 5597 -912 12229 -907
rect 5597 -1008 5799 -912
rect 6326 -999 12229 -912
rect 6326 -1008 6343 -999
rect 5597 -1019 6343 -1008
rect 5597 -1021 5776 -1019
rect 6272 -1021 6343 -1019
rect 5612 -1906 6906 -1863
rect 5612 -1940 5800 -1906
rect 6838 -1940 6906 -1906
rect 5612 -1948 6906 -1940
rect 5612 -1966 5812 -1948
rect 5612 -2324 5740 -1966
rect 5774 -2324 5812 -1966
rect 5612 -2341 5812 -2324
rect 6825 -1966 6906 -1948
rect 6825 -2324 6864 -1966
rect 6898 -2324 6906 -1966
rect 6825 -2341 6906 -2324
rect 5612 -2350 6906 -2341
rect 5612 -2384 5800 -2350
rect 6838 -2384 6906 -2350
rect 5612 -2426 6906 -2384
rect 5612 -2555 7151 -2426
rect 5612 -2556 6545 -2555
rect 5612 -2696 5648 -2556
rect 6726 -2695 7151 -2555
rect 6550 -2696 7151 -2695
rect 5612 -2751 7151 -2696
<< viali >>
rect 5614 2053 12192 2190
rect 5614 2019 5690 2053
rect 5690 2019 12146 2053
rect 12146 2019 12192 2053
rect 5614 2016 12192 2019
rect 5807 -776 12146 -751
rect 12146 -776 12148 -751
rect 5807 -863 12148 -776
rect 5799 -1008 6326 -912
rect 6545 -2556 6726 -2555
rect 5648 -2695 6726 -2556
rect 5648 -2696 6550 -2695
<< metal1 >>
rect 5602 2190 12204 2196
rect 5602 2016 5614 2190
rect 12192 2016 12204 2190
rect 5602 2010 12204 2016
rect 5811 1565 5821 1765
rect 5885 1565 5895 1765
rect 5935 943 6024 1812
rect 6074 1809 6164 1855
rect 6073 989 6083 1189
rect 6139 989 6149 1189
rect 6199 948 6288 1810
rect 6448 1413 6537 1812
rect 6589 1809 6665 1855
rect 6591 1565 6601 1765
rect 6653 1565 6663 1765
rect 6333 1313 6343 1413
rect 6395 1313 6405 1413
rect 6448 1313 6467 1413
rect 6519 1313 6537 1413
rect 6077 899 6147 945
rect 6199 941 6224 948
rect 6214 896 6224 941
rect 6324 896 6334 948
rect 6448 943 6537 1313
rect 6712 1413 6800 1816
rect 6712 1313 6732 1413
rect 6784 1313 6800 1413
rect 6849 1313 6859 1413
rect 6911 1313 6921 1413
rect 6712 948 6800 1313
rect 6591 899 6681 945
rect 6712 939 6740 948
rect 6730 896 6740 939
rect 6840 896 6850 948
rect 6973 939 7061 1816
rect 7105 1809 7182 1855
rect 7105 989 7115 1189
rect 7171 989 7181 1189
rect 7107 899 7184 945
rect 7236 943 7324 1820
rect 7365 1809 7439 1855
rect 7359 1565 7369 1765
rect 7433 1565 7443 1765
rect 7365 899 7439 945
rect 7486 941 7574 1818
rect 7624 1809 7703 1855
rect 7621 989 7631 1189
rect 7687 989 7697 1189
rect 7745 958 7833 1820
rect 7998 1414 8091 1815
rect 8140 1809 8213 1855
rect 8139 1565 8149 1765
rect 8201 1565 8211 1765
rect 7881 1313 7891 1413
rect 7943 1313 7953 1413
rect 7998 1314 8014 1414
rect 8066 1314 8091 1414
rect 7723 948 7833 958
rect 7625 899 7714 945
rect 7723 896 7746 948
rect 7872 896 7882 948
rect 7998 941 8091 1314
rect 8260 1412 8348 1816
rect 8260 1312 8276 1412
rect 8328 1312 8348 1412
rect 8397 1313 8407 1413
rect 8459 1313 8469 1413
rect 8260 948 8348 1312
rect 8140 899 8213 945
rect 8260 939 8288 948
rect 8278 896 8288 939
rect 8388 896 8398 948
rect 8525 943 8613 1820
rect 8655 1809 8728 1855
rect 8653 989 8663 1189
rect 8719 989 8729 1189
rect 8655 899 8728 945
rect 8781 941 8869 1818
rect 8915 1809 8988 1855
rect 8907 1565 8917 1765
rect 8981 1565 8991 1765
rect 8915 899 8988 945
rect 9038 943 9126 1820
rect 9170 1809 9242 1855
rect 9169 989 9179 1189
rect 9235 989 9245 1189
rect 9297 948 9385 1820
rect 9429 1313 9439 1413
rect 9491 1313 9501 1413
rect 9549 1411 9637 1816
rect 9688 1809 9760 1855
rect 9686 1565 9696 1765
rect 9748 1565 9758 1765
rect 9549 1311 9569 1411
rect 9621 1311 9637 1411
rect 9172 899 9263 945
rect 9280 896 9294 948
rect 9420 896 9430 948
rect 9549 939 9637 1311
rect 9806 1414 9894 1818
rect 9806 1314 9821 1414
rect 9873 1314 9894 1414
rect 9806 948 9894 1314
rect 9945 1313 9955 1413
rect 10007 1313 10017 1413
rect 9688 899 9760 945
rect 9806 941 9836 948
rect 9826 896 9836 941
rect 9936 896 9946 948
rect 10073 941 10161 1818
rect 10205 1809 10277 1855
rect 10201 989 10211 1189
rect 10267 989 10277 1189
rect 10205 899 10277 945
rect 10317 941 10405 1818
rect 10462 1809 10533 1855
rect 10455 1565 10465 1765
rect 10529 1565 10539 1765
rect 10462 899 10533 945
rect 10582 941 10670 1818
rect 10720 1809 10793 1855
rect 10732 1285 10778 1441
rect 10717 989 10727 1189
rect 10783 989 10793 1189
rect 10833 948 10921 1820
rect 11099 1416 11187 1820
rect 11237 1809 11307 1855
rect 11235 1565 11245 1765
rect 11297 1565 11307 1765
rect 10977 1313 10987 1413
rect 11039 1313 11049 1413
rect 11099 1316 11112 1416
rect 11164 1316 11187 1416
rect 10990 977 11036 1255
rect 10720 899 10800 945
rect 10833 943 10843 948
rect 10837 896 10843 943
rect 10968 945 10978 948
rect 10968 899 10980 945
rect 11046 899 11049 945
rect 11099 943 11187 1316
rect 11356 1419 11444 1822
rect 11356 1314 11374 1419
rect 11426 1314 11444 1419
rect 11356 948 11444 1314
rect 11493 1313 11503 1413
rect 11555 1313 11565 1413
rect 11356 945 11384 948
rect 11237 899 11307 945
rect 10968 896 10978 899
rect 11374 896 11384 945
rect 11484 896 11494 948
rect 11630 941 11718 1818
rect 11752 1809 11823 1855
rect 11749 989 11759 1189
rect 11815 989 11825 1189
rect 11873 948 11961 1818
rect 12003 1565 12013 1765
rect 12077 1565 12087 1765
rect 11752 899 11823 945
rect 11873 941 11900 948
rect 11890 896 11900 941
rect 12000 896 12010 948
rect 7723 886 7768 896
rect 5701 670 6272 722
rect 6372 670 7046 722
rect 7146 670 7820 722
rect 7920 670 8594 722
rect 8694 670 9368 722
rect 9468 670 10142 722
rect 10242 670 10916 722
rect 11016 670 11690 722
rect 11790 670 11948 722
rect 12048 670 12058 722
rect 5701 -1470 5753 670
rect 5892 525 6014 577
rect 6114 525 6788 577
rect 6888 525 7562 577
rect 7662 525 8336 577
rect 8436 525 9110 577
rect 9210 525 9884 577
rect 9984 525 10658 577
rect 10758 525 11432 577
rect 11532 525 11948 577
rect 12048 525 12058 577
rect 5956 336 5966 377
rect 5943 325 5966 336
rect 6066 325 6076 377
rect 6888 374 6898 377
rect 5943 -19 6031 325
rect 5943 -119 5962 -19
rect 6014 -119 6031 -19
rect 6075 -117 6085 -17
rect 6137 -117 6147 -17
rect 5817 -492 5827 -292
rect 5879 -492 5889 -292
rect 5943 -541 6031 -119
rect 6195 -539 6283 338
rect 6334 328 6403 374
rect 6331 -491 6341 -291
rect 6397 -491 6407 -291
rect 6335 -582 6404 -536
rect 6444 -541 6532 336
rect 6593 328 6662 374
rect 6585 84 6595 284
rect 6659 84 6669 284
rect 6589 -582 6663 -536
rect 6714 -539 6802 338
rect 6850 328 6898 374
rect 6888 325 6898 328
rect 7098 325 7108 377
rect 6847 -492 6857 -292
rect 6913 -492 6923 -292
rect 6850 -582 6922 -536
rect 6963 -537 7051 325
rect 7226 -16 7314 338
rect 7366 328 7436 374
rect 7504 336 7514 377
rect 7107 -117 7117 -17
rect 7169 -117 7179 -17
rect 7226 -116 7240 -16
rect 7292 -116 7314 -16
rect 7226 -539 7314 -116
rect 7480 325 7514 336
rect 7614 325 7624 377
rect 8452 374 8462 377
rect 7480 -15 7568 325
rect 7480 -115 7496 -15
rect 7548 -115 7568 -15
rect 7365 -492 7375 -292
rect 7427 -492 7437 -292
rect 7366 -582 7436 -536
rect 7480 -541 7568 -115
rect 7623 -117 7633 -17
rect 7685 -117 7695 -17
rect 7747 -541 7835 336
rect 7882 328 7952 374
rect 7879 -492 7889 -292
rect 7945 -492 7955 -292
rect 7881 -582 7951 -536
rect 8000 -539 8088 338
rect 8141 328 8211 374
rect 8133 84 8143 284
rect 8207 84 8217 284
rect 8140 -582 8210 -536
rect 8252 -539 8340 338
rect 8399 328 8462 374
rect 8452 325 8462 328
rect 8646 325 8656 377
rect 8395 -492 8405 -292
rect 8461 -492 8471 -292
rect 8399 -582 8468 -536
rect 8523 -541 8611 325
rect 8769 -17 8850 333
rect 8913 328 8985 374
rect 9052 331 9062 377
rect 8655 -117 8665 -17
rect 8717 -117 8727 -17
rect 8769 -117 8782 -17
rect 8834 -117 8850 -17
rect 8769 -541 8850 -117
rect 9029 325 9062 331
rect 9162 325 9172 377
rect 10000 374 10010 377
rect 9029 -19 9110 325
rect 9029 -119 9044 -19
rect 9096 -119 9110 -19
rect 9171 -116 9181 -16
rect 9233 -116 9243 -16
rect 8913 -492 8923 -292
rect 8975 -492 8985 -292
rect 8914 -582 8986 -536
rect 9029 -543 9110 -119
rect 9291 -539 9379 338
rect 9430 328 9523 374
rect 9427 -492 9437 -292
rect 9493 -492 9503 -292
rect 9431 -582 9502 -536
rect 9547 -539 9635 338
rect 9678 328 9760 374
rect 9681 84 9691 284
rect 9755 84 9765 284
rect 9687 -582 9760 -536
rect 9808 -539 9896 338
rect 9947 328 10010 374
rect 10000 325 10010 328
rect 10194 325 10204 377
rect 9943 -492 9953 -292
rect 10009 -492 10019 -292
rect 9945 -582 10017 -536
rect 10063 -539 10151 325
rect 10203 -117 10213 -17
rect 10265 -117 10275 -17
rect 10318 -19 10424 337
rect 10463 328 10534 374
rect 10600 334 10610 377
rect 10318 -119 10340 -19
rect 10392 -119 10424 -19
rect 10318 -539 10424 -119
rect 10573 325 10610 334
rect 10710 325 10720 377
rect 11548 374 11558 377
rect 10573 -17 10679 325
rect 10573 -117 10595 -17
rect 10647 -117 10679 -17
rect 10719 -117 10729 -17
rect 10781 -117 10791 -17
rect 10461 -492 10471 -292
rect 10523 -492 10533 -292
rect 10461 -582 10532 -536
rect 10573 -542 10679 -117
rect 10843 -539 10931 338
rect 10977 328 11046 374
rect 10975 -492 10985 -292
rect 11041 -492 11051 -292
rect 10979 -582 11048 -536
rect 11099 -541 11187 336
rect 11235 328 11307 374
rect 11229 84 11239 284
rect 11303 84 11313 284
rect 11236 -582 11308 -536
rect 11358 -539 11446 338
rect 11494 328 11558 374
rect 11548 325 11558 328
rect 11742 325 11752 377
rect 11890 336 11900 377
rect 11871 325 11900 336
rect 12000 325 12010 377
rect 11491 -492 11501 -292
rect 11557 -492 11567 -292
rect 11495 -582 11564 -536
rect 11618 -541 11706 325
rect 11871 -15 11959 325
rect 11751 -117 11761 -17
rect 11813 -117 11823 -17
rect 11871 -115 11887 -15
rect 11939 -115 11959 -15
rect 11871 -541 11959 -115
rect 12009 -492 12019 -292
rect 12071 -492 12081 -292
rect 5794 -751 12160 -745
rect 5794 -863 5807 -751
rect 12148 -863 12160 -751
rect 5794 -869 12160 -863
rect 5787 -912 6338 -906
rect 5787 -1008 5799 -912
rect 6326 -1008 6338 -912
rect 5787 -1014 6338 -1008
rect 5701 -1522 5915 -1470
rect 5905 -1584 5915 -1522
rect 5967 -1522 6178 -1470
rect 5967 -1584 5977 -1522
rect 6039 -2045 6049 -1984
rect 6016 -2050 6049 -2045
rect 6643 -2050 6653 -1984
rect 5905 -2185 5915 -2109
rect 5967 -2185 5977 -2109
rect 6016 -2246 6120 -2050
rect 6162 -2056 6236 -2050
rect 6163 -2185 6173 -2109
rect 6225 -2185 6235 -2109
rect 6165 -2284 6235 -2238
rect 6271 -2244 6375 -2050
rect 6423 -2056 6497 -2050
rect 6434 -2238 6480 -2056
rect 6423 -2284 6493 -2238
rect 6539 -2246 6643 -2050
rect 6681 -2056 6917 -2010
rect 6679 -2185 6689 -2109
rect 6741 -2185 6751 -2109
rect 6533 -2550 6738 -2549
rect 5636 -2555 6738 -2550
rect 5636 -2556 6545 -2555
rect 5636 -2696 5648 -2556
rect 6726 -2695 6738 -2555
rect 6550 -2696 6738 -2695
rect 5636 -2701 6738 -2696
rect 5636 -2702 6562 -2701
<< via1 >>
rect 5614 2016 12192 2190
rect 5821 1565 5885 1765
rect 6083 989 6139 1189
rect 6601 1565 6653 1765
rect 6343 1313 6395 1413
rect 6467 1313 6519 1413
rect 6224 896 6324 948
rect 6732 1313 6784 1413
rect 6859 1313 6911 1413
rect 6740 896 6840 948
rect 7115 989 7171 1189
rect 7369 1565 7433 1765
rect 7631 989 7687 1189
rect 8149 1565 8201 1765
rect 7891 1313 7943 1413
rect 8014 1314 8066 1414
rect 7746 896 7872 948
rect 8276 1312 8328 1412
rect 8407 1313 8459 1413
rect 8288 896 8388 948
rect 8663 989 8719 1189
rect 8917 1565 8981 1765
rect 9179 989 9235 1189
rect 9439 1313 9491 1413
rect 9696 1565 9748 1765
rect 9569 1311 9621 1411
rect 9294 896 9420 948
rect 9821 1314 9873 1414
rect 9955 1313 10007 1413
rect 9836 896 9936 948
rect 10211 989 10267 1189
rect 10465 1565 10529 1765
rect 10727 989 10783 1189
rect 11245 1565 11297 1765
rect 10987 1313 11039 1413
rect 11112 1316 11164 1416
rect 10843 896 10968 948
rect 11374 1314 11426 1419
rect 11503 1313 11555 1413
rect 11384 896 11484 948
rect 11759 989 11815 1189
rect 12013 1565 12077 1765
rect 11900 896 12000 948
rect 6272 670 6372 722
rect 7046 670 7146 722
rect 7820 670 7920 722
rect 8594 670 8694 722
rect 9368 670 9468 722
rect 10142 670 10242 722
rect 10916 670 11016 722
rect 11690 670 11790 722
rect 11948 670 12048 722
rect 6014 525 6114 577
rect 6788 525 6888 577
rect 7562 525 7662 577
rect 8336 525 8436 577
rect 9110 525 9210 577
rect 9884 525 9984 577
rect 10658 525 10758 577
rect 11432 525 11532 577
rect 11948 525 12048 577
rect 5966 325 6066 377
rect 5962 -119 6014 -19
rect 6085 -117 6137 -17
rect 5827 -492 5879 -292
rect 6341 -491 6397 -291
rect 6595 84 6659 284
rect 6898 325 7098 377
rect 6857 -492 6913 -292
rect 7117 -117 7169 -17
rect 7240 -116 7292 -16
rect 7514 325 7614 377
rect 7496 -115 7548 -15
rect 7375 -492 7427 -292
rect 7633 -117 7685 -17
rect 7889 -492 7945 -292
rect 8143 84 8207 284
rect 8462 325 8646 377
rect 8405 -492 8461 -292
rect 8665 -117 8717 -17
rect 8782 -117 8834 -17
rect 9062 325 9162 377
rect 9044 -119 9096 -19
rect 9181 -116 9233 -16
rect 8923 -492 8975 -292
rect 9437 -492 9493 -292
rect 9691 84 9755 284
rect 10010 325 10194 377
rect 9953 -492 10009 -292
rect 10213 -117 10265 -17
rect 10340 -119 10392 -19
rect 10610 325 10710 377
rect 10595 -117 10647 -17
rect 10729 -117 10781 -17
rect 10471 -492 10523 -292
rect 10985 -492 11041 -292
rect 11239 84 11303 284
rect 11558 325 11742 377
rect 11900 325 12000 377
rect 11501 -492 11557 -292
rect 11761 -117 11813 -17
rect 11887 -115 11939 -15
rect 12019 -492 12071 -292
rect 5807 -863 12148 -751
rect 5799 -1008 6326 -912
rect 5915 -1584 5967 -1470
rect 6049 -2050 6643 -1984
rect 5915 -2185 5967 -2109
rect 6173 -2185 6225 -2109
rect 6689 -2185 6741 -2109
rect 6545 -2556 6726 -2555
rect 5648 -2695 6726 -2556
rect 5648 -2696 6550 -2695
<< metal2 >>
rect 5511 2190 12192 2200
rect 5511 2016 5614 2190
rect 5511 2006 12192 2016
rect 5821 1765 5885 1775
rect 5821 1555 5885 1565
rect 6601 1765 6653 2006
rect 6601 1555 6653 1565
rect 7369 1765 7433 1775
rect 7369 1555 7433 1565
rect 8149 1765 8201 2006
rect 8149 1555 8201 1565
rect 8917 1765 8981 1775
rect 8917 1555 8981 1565
rect 9696 1765 9748 2006
rect 9696 1555 9748 1565
rect 10465 1765 10529 1775
rect 10465 1555 10529 1565
rect 11245 1765 11297 2006
rect 11245 1555 11297 1565
rect 12013 1765 12077 1775
rect 12013 1555 12077 1565
rect 8014 1423 8066 1424
rect 9821 1423 9873 1424
rect 11112 1423 11164 1426
rect 11374 1423 11426 1424
rect 6343 1419 12351 1423
rect 6343 1416 11374 1419
rect 6343 1414 11112 1416
rect 6343 1413 8014 1414
rect 6395 1313 6467 1413
rect 6519 1313 6732 1413
rect 6784 1313 6859 1413
rect 6911 1313 7891 1413
rect 7943 1314 8014 1413
rect 8066 1413 9821 1414
rect 8066 1412 8407 1413
rect 8066 1314 8276 1412
rect 7943 1313 8276 1314
rect 6343 1312 8276 1313
rect 8328 1313 8407 1412
rect 8459 1313 9439 1413
rect 9491 1411 9821 1413
rect 9491 1313 9569 1411
rect 8328 1312 9569 1313
rect 6343 1311 9569 1312
rect 9621 1314 9821 1411
rect 9873 1413 11112 1414
rect 9873 1314 9955 1413
rect 9621 1313 9955 1314
rect 10007 1313 10987 1413
rect 11039 1316 11112 1413
rect 11164 1316 11374 1416
rect 11039 1314 11374 1316
rect 11426 1413 12351 1419
rect 11426 1314 11503 1413
rect 11039 1313 11503 1314
rect 11555 1313 12351 1413
rect 9621 1311 12351 1313
rect 6343 1303 12351 1311
rect 8276 1302 8328 1303
rect 9569 1301 9621 1303
rect 6083 1189 6139 1199
rect 6083 979 6139 989
rect 7115 1189 7171 1199
rect 7115 979 7171 989
rect 7631 1189 7687 1199
rect 7631 979 7687 989
rect 8663 1189 8719 1199
rect 8663 979 8719 989
rect 9179 1189 9235 1199
rect 9179 979 9235 989
rect 10211 1189 10267 1199
rect 10211 979 10267 989
rect 10727 1189 10783 1199
rect 10727 979 10783 989
rect 11759 1189 11815 1199
rect 11759 979 11815 989
rect 6224 948 6324 958
rect 6224 886 6324 896
rect 6740 948 6840 958
rect 6740 886 6840 896
rect 7740 948 7872 958
rect 7740 896 7746 948
rect 7740 886 7872 896
rect 8288 948 8388 958
rect 8288 886 8388 896
rect 9294 948 9420 958
rect 9294 886 9420 896
rect 9836 948 9936 958
rect 9836 886 9936 896
rect 10843 948 10968 958
rect 10843 886 10968 896
rect 11384 948 11484 958
rect 11384 886 11484 896
rect 11900 948 12000 958
rect 11900 886 12000 896
rect 6272 732 6324 886
rect 6272 722 6372 732
rect 6272 660 6372 670
rect 6788 587 6840 886
rect 7820 732 7872 886
rect 7046 722 7146 732
rect 7046 660 7146 670
rect 7820 722 7920 732
rect 7820 660 7920 670
rect 6014 577 6114 587
rect 6014 515 6114 525
rect 6788 577 6888 587
rect 6788 515 6888 525
rect 6014 387 6066 515
rect 7046 387 7098 660
rect 8336 587 8388 886
rect 9368 732 9420 886
rect 8594 722 8694 732
rect 8594 660 8694 670
rect 9368 722 9468 732
rect 9368 660 9468 670
rect 7562 577 7662 587
rect 7562 515 7662 525
rect 8336 577 8436 587
rect 8336 515 8436 525
rect 7562 387 7614 515
rect 8594 387 8646 660
rect 9884 587 9936 886
rect 10916 732 10968 886
rect 10142 722 10242 732
rect 10142 660 10242 670
rect 10916 722 11016 732
rect 10916 660 11016 670
rect 9110 577 9210 587
rect 9110 515 9210 525
rect 9884 577 9984 587
rect 9884 515 9984 525
rect 9110 387 9162 515
rect 10142 387 10194 660
rect 11432 587 11484 886
rect 11948 732 12000 886
rect 11690 722 11790 732
rect 11690 660 11790 670
rect 11948 722 12048 732
rect 11948 660 12048 670
rect 10658 577 10758 587
rect 10658 515 10758 525
rect 11432 577 11532 587
rect 11432 515 11532 525
rect 10658 387 10710 515
rect 11690 387 11742 660
rect 11948 577 12048 587
rect 11948 515 12048 525
rect 11948 387 12000 515
rect 5966 377 6066 387
rect 5966 315 6066 325
rect 6898 377 7098 387
rect 6898 315 7098 325
rect 7514 377 7614 387
rect 7514 315 7614 325
rect 8462 377 8646 387
rect 8462 315 8646 325
rect 9062 377 9162 387
rect 9062 315 9162 325
rect 10010 377 10194 387
rect 10010 315 10194 325
rect 10610 377 10710 387
rect 10610 315 10710 325
rect 11558 377 11742 387
rect 11558 315 11742 325
rect 11900 377 12000 387
rect 11900 315 12000 325
rect 6595 284 6659 294
rect 6595 74 6659 84
rect 8143 284 8207 294
rect 8143 74 8207 84
rect 9691 284 9755 294
rect 9691 74 9755 84
rect 11239 284 11303 294
rect 11239 74 11303 84
rect 7240 -7 7292 -6
rect 7496 -7 7548 -5
rect 9181 -7 9233 -6
rect 11887 -7 11939 -5
rect 12231 -7 12351 1303
rect 5938 -15 12351 -7
rect 5938 -16 7496 -15
rect 5938 -17 7240 -16
rect 5938 -19 6085 -17
rect 5938 -119 5962 -19
rect 6014 -117 6085 -19
rect 6137 -117 7117 -17
rect 7169 -116 7240 -17
rect 7292 -115 7496 -16
rect 7548 -16 11887 -15
rect 7548 -17 9181 -16
rect 7548 -115 7633 -17
rect 7292 -116 7633 -115
rect 7169 -117 7633 -116
rect 7685 -117 8665 -17
rect 8717 -117 8782 -17
rect 8834 -19 9181 -17
rect 8834 -117 9044 -19
rect 6014 -119 9044 -117
rect 9096 -116 9181 -19
rect 9233 -17 11887 -16
rect 9233 -116 10213 -17
rect 9096 -117 10213 -116
rect 10265 -19 10595 -17
rect 10265 -117 10340 -19
rect 9096 -119 10340 -117
rect 10392 -117 10595 -19
rect 10647 -117 10729 -17
rect 10781 -117 11761 -17
rect 11813 -115 11887 -17
rect 11939 -115 12351 -15
rect 11813 -117 12351 -115
rect 10392 -119 12351 -117
rect 5938 -127 12351 -119
rect 5962 -129 6014 -127
rect 9044 -129 9096 -127
rect 10340 -129 10392 -127
rect 5827 -292 5879 -282
rect 5827 -741 5879 -492
rect 6341 -291 6397 -281
rect 6341 -501 6397 -491
rect 6857 -292 6913 -282
rect 6857 -502 6913 -492
rect 7375 -292 7427 -282
rect 7375 -741 7427 -492
rect 7889 -292 7945 -282
rect 7889 -502 7945 -492
rect 8405 -292 8461 -282
rect 8405 -502 8461 -492
rect 8923 -292 8975 -282
rect 8923 -741 8975 -492
rect 9437 -292 9493 -282
rect 9437 -502 9493 -492
rect 9953 -292 10009 -282
rect 9953 -502 10009 -492
rect 10471 -292 10523 -282
rect 10471 -741 10523 -492
rect 10985 -292 11041 -282
rect 10985 -502 11041 -492
rect 11501 -292 11557 -282
rect 11501 -502 11557 -492
rect 12019 -292 12071 -282
rect 12019 -741 12071 -492
rect 5794 -751 12148 -741
rect 5794 -863 5807 -751
rect 5794 -873 12148 -863
rect 5794 -912 6326 -873
rect 5794 -1008 5799 -912
rect 5794 -1018 6326 -1008
rect 6395 -1236 6457 -1235
rect 6389 -1245 6465 -1236
rect 6389 -1364 6395 -1245
rect 6457 -1312 6465 -1245
rect 6457 -1364 6497 -1312
rect 6389 -1392 6497 -1364
rect 5915 -1470 5967 -1460
rect 5915 -2109 5967 -1584
rect 6049 -1984 6643 -1974
rect 6049 -2060 6643 -2050
rect 5915 -2195 5967 -2185
rect 6173 -2109 6225 -2099
rect 6173 -2546 6225 -2185
rect 6689 -2109 6741 -2099
rect 6689 -2545 6741 -2185
rect 6545 -2546 6741 -2545
rect 5613 -2555 6741 -2546
rect 5613 -2556 6545 -2555
rect 5613 -2696 5648 -2556
rect 6726 -2695 6741 -2555
rect 6550 -2696 6741 -2695
rect 5613 -2705 6741 -2696
rect 5613 -2706 6550 -2705
<< via2 >>
rect 5821 1565 5885 1765
rect 7369 1565 7433 1765
rect 8917 1565 8981 1765
rect 10465 1565 10529 1765
rect 12013 1565 12077 1765
rect 6083 989 6139 1189
rect 7115 989 7171 1189
rect 7631 989 7687 1189
rect 8663 989 8719 1189
rect 9179 989 9235 1189
rect 10211 989 10267 1189
rect 10727 989 10783 1189
rect 11759 989 11815 1189
rect 6595 84 6659 284
rect 8143 84 8207 284
rect 9691 84 9755 284
rect 11239 84 11303 284
rect 6341 -491 6397 -291
rect 6857 -492 6913 -292
rect 7889 -492 7945 -292
rect 8405 -492 8461 -292
rect 9437 -492 9493 -292
rect 9953 -492 10009 -292
rect 10985 -492 11041 -292
rect 11501 -492 11557 -292
rect 6395 -1364 6457 -1245
rect 6049 -2050 6643 -1984
<< metal3 >>
rect 5811 1765 5895 1770
rect 5811 1565 5821 1765
rect 5885 1565 5895 1765
rect 5811 1560 5895 1565
rect 7359 1765 7443 1770
rect 7359 1565 7369 1765
rect 7433 1565 7443 1765
rect 7359 1560 7443 1565
rect 8907 1765 8991 1770
rect 8907 1565 8917 1765
rect 8981 1565 8991 1765
rect 8907 1560 8991 1565
rect 10455 1765 10539 1770
rect 10455 1565 10465 1765
rect 10529 1565 10539 1765
rect 10455 1560 10539 1565
rect 12003 1765 12087 1770
rect 12003 1565 12013 1765
rect 12077 1565 12087 1765
rect 12003 1560 12087 1565
rect 6073 1189 6149 1194
rect 6073 1060 6083 1189
rect 5683 989 6083 1060
rect 6139 1060 6149 1189
rect 7105 1189 7181 1194
rect 7105 1060 7115 1189
rect 6139 989 7115 1060
rect 7171 1060 7181 1189
rect 7621 1189 7697 1194
rect 7621 1060 7631 1189
rect 7171 989 7631 1060
rect 7687 1060 7697 1189
rect 8653 1189 8729 1194
rect 8653 1060 8663 1189
rect 7687 989 8663 1060
rect 8719 1060 8729 1189
rect 9169 1189 9245 1194
rect 9169 1060 9179 1189
rect 8719 989 9179 1060
rect 9235 1060 9245 1189
rect 10201 1189 10277 1194
rect 10201 1060 10211 1189
rect 9235 989 10211 1060
rect 10267 1060 10277 1189
rect 10717 1189 10793 1194
rect 10717 1060 10727 1189
rect 10267 989 10727 1060
rect 10783 1060 10793 1189
rect 11749 1189 11825 1194
rect 11749 1060 11759 1189
rect 10783 989 11759 1060
rect 11815 989 11825 1189
rect 5683 986 11825 989
rect 5683 -421 5757 986
rect 6073 984 6149 986
rect 7105 984 7181 986
rect 7621 984 7697 986
rect 8653 984 8729 986
rect 9169 984 9245 986
rect 10201 984 10277 986
rect 10717 984 10793 986
rect 11685 984 11825 986
rect 6585 284 6669 289
rect 6585 84 6595 284
rect 6659 84 6669 284
rect 6585 79 6669 84
rect 8133 284 8217 289
rect 8133 84 8143 284
rect 8207 84 8217 284
rect 8133 79 8217 84
rect 9681 284 9765 289
rect 9681 84 9691 284
rect 9755 84 9765 284
rect 9681 79 9765 84
rect 11229 284 11313 289
rect 11229 84 11239 284
rect 11303 84 11313 284
rect 11229 79 11313 84
rect 6331 -291 6407 -286
rect 6331 -421 6341 -291
rect 5683 -491 6341 -421
rect 6397 -421 6407 -291
rect 6847 -292 6923 -287
rect 6847 -421 6857 -292
rect 6397 -491 6857 -421
rect 5683 -492 6857 -491
rect 6913 -421 6923 -292
rect 7879 -292 7955 -287
rect 7879 -421 7889 -292
rect 6913 -492 7889 -421
rect 7945 -421 7955 -292
rect 8395 -292 8471 -287
rect 8395 -421 8405 -292
rect 7945 -492 8405 -421
rect 8461 -421 8471 -292
rect 9427 -292 9503 -287
rect 9427 -421 9437 -292
rect 8461 -492 9437 -421
rect 9493 -421 9503 -292
rect 9943 -292 10019 -287
rect 9943 -421 9953 -292
rect 9493 -492 9953 -421
rect 10009 -421 10019 -292
rect 10975 -292 11051 -287
rect 10975 -421 10985 -292
rect 10009 -492 10985 -421
rect 11041 -421 11051 -292
rect 11491 -292 11567 -287
rect 11491 -421 11501 -292
rect 11041 -492 11501 -421
rect 11557 -492 11567 -292
rect 5683 -497 11567 -492
rect 6385 -1245 6467 -497
rect 6385 -1364 6395 -1245
rect 6457 -1364 6467 -1245
rect 6385 -1369 6467 -1364
rect 6039 -1984 6653 -1979
rect 6039 -2050 6049 -1984
rect 6643 -2050 6653 -1984
rect 6039 -2055 6653 -2050
<< via3 >>
rect 5821 1565 5885 1765
rect 7369 1565 7433 1765
rect 8917 1565 8981 1765
rect 10465 1565 10529 1765
rect 12013 1565 12077 1765
rect 6595 84 6659 284
rect 8143 84 8207 284
rect 9691 84 9755 284
rect 11239 84 11303 284
rect 6049 -2050 6643 -1984
<< metal4 >>
rect 5537 1765 12078 1766
rect 5537 1690 5821 1765
rect 5537 1035 5613 1690
rect 5820 1565 5821 1690
rect 5885 1690 7369 1765
rect 5885 1565 5886 1690
rect 5820 1564 5886 1565
rect 7368 1565 7369 1690
rect 7433 1690 8917 1765
rect 7433 1565 7434 1690
rect 7368 1564 7434 1565
rect 8916 1565 8917 1690
rect 8981 1690 10465 1765
rect 8981 1565 8982 1690
rect 8916 1564 8982 1565
rect 10464 1565 10465 1690
rect 10529 1690 12013 1765
rect 10529 1565 10530 1690
rect 10464 1564 10530 1565
rect 12012 1565 12013 1690
rect 12077 1565 12078 1765
rect 12012 1564 12078 1565
rect 5349 958 5613 1035
rect 5349 -1980 5425 958
rect 5537 285 5613 958
rect 5537 284 11304 285
rect 5537 209 6595 284
rect 6594 84 6595 209
rect 6659 209 8143 284
rect 6659 84 6660 209
rect 6594 83 6660 84
rect 8142 84 8143 209
rect 8207 209 9691 284
rect 8207 84 8208 209
rect 8142 83 8208 84
rect 9690 84 9691 209
rect 9755 209 11239 284
rect 9755 84 9756 209
rect 9690 83 9756 84
rect 11238 84 11239 209
rect 11303 84 11304 284
rect 11238 83 11304 84
rect 5349 -1984 6670 -1980
rect 5349 -2050 6049 -1984
rect 6643 -2050 6670 -1984
rect 5349 -2056 6670 -2050
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2_0 ~/Dalin/Projects/tinytape/voltage_ref/stge -1 backup1/layout_stage-1
timestamp 1738283136
transform 1 0 11916 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__pfet_01v8_lvt_SCQJZQ  sky130_fd_pr__pfet_01v8_lvt_SCQJZQ_0 ~/Dalin/Projects/tinytape/voltage_ref/stge -1 backup1/layout_stage-1
timestamp 1738536365
transform 1 0 6586 0 1 -2147
box -194 -150 194 150
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM1
timestamp 1738283136
transform 1 0 6498 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM2
timestamp 1738283136
transform 1 0 6240 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM3
timestamp 1738283136
transform 1 0 5982 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM4
timestamp 1738283136
transform 1 0 7272 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM5
timestamp 1738283136
transform 1 0 7530 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM6
timestamp 1738283136
transform 1 0 8820 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM7
timestamp 1738283136
transform 1 0 9078 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__pfet_01v8_lvt_SCQJZQ  XM8
timestamp 1738536365
transform 1 0 6328 0 1 -2147
box -194 -150 194 150
use sky130_fd_pr__pfet_01v8_lvt_SCQJZQ  XM9
timestamp 1738536365
transform 1 0 6070 0 1 -2147
box -194 -150 194 150
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM10
timestamp 1738283136
transform 1 0 10368 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM11
timestamp 1738283136
transform 1 0 10626 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM12
timestamp 1738283136
transform 1 0 11916 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM14
timestamp 1738283136
transform 1 0 6498 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM15
timestamp 1738283136
transform 1 0 6756 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM16
timestamp 1738283136
transform 1 0 8046 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM17
timestamp 1738283136
transform 1 0 8304 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM18
timestamp 1738283136
transform 1 0 9594 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM19
timestamp 1738283136
transform 1 0 9852 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM20
timestamp 1738283136
transform 1 0 11142 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM21
timestamp 1738283136
transform 1 0 11400 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM22
timestamp 1738283136
transform 1 0 7014 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM23
timestamp 1738283136
transform 1 0 7788 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM24
timestamp 1738283136
transform 1 0 8562 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM25
timestamp 1738283136
transform 1 0 9336 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM26
timestamp 1738283136
transform 1 0 10110 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM27
timestamp 1738283136
transform 1 0 10884 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM28
timestamp 1738283136
transform 1 0 11658 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM29
timestamp 1738283136
transform 1 0 6240 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM30
timestamp 1738283136
transform 1 0 7014 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM31
timestamp 1738283136
transform 1 0 7788 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM32
timestamp 1738283136
transform 1 0 8562 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM33
timestamp 1738283136
transform 1 0 9336 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM34
timestamp 1738283136
transform 1 0 10110 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM35
timestamp 1738283136
transform 1 0 10884 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM36
timestamp 1738283136
transform 1 0 6756 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM37
timestamp 1738283136
transform 1 0 8046 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM38
timestamp 1738283136
transform 1 0 8304 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM39
timestamp 1738283136
transform 1 0 9594 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM40
timestamp 1738283136
transform 1 0 9852 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM41
timestamp 1738283136
transform 1 0 11142 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM42
timestamp 1738283136
transform 1 0 11400 0 1 1377
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM43
timestamp 1738283136
transform 1 0 5982 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM44
timestamp 1738283136
transform 1 0 7272 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM45
timestamp 1738283136
transform 1 0 7530 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM46
timestamp 1738283136
transform 1 0 8820 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM47
timestamp 1738283136
transform 1 0 9078 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM48
timestamp 1738283136
transform 1 0 10368 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM49
timestamp 1738283136
transform 1 0 10626 0 1 -104
box -158 -488 158 488
use sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2  XM50
timestamp 1738283136
transform 1 0 11658 0 1 -104
box -158 -488 158 488
<< labels >>
rlabel metal2 5614 -2623 5614 -2623 3 vcc
port 1 e
rlabel metal2 5512 2112 5512 2112 3 vss
port 2 e
rlabel metal2 6496 -1351 6496 -1351 3 vref0
port 3 e
rlabel metal1 6916 -2033 6916 -2033 3 vr
port 4 e
rlabel metal1 6176 -1495 6176 -1495 3 vd
port 5 e
<< end >>
