* NGSPICE file created from 3rd_3_OTA_flat.ext - technology: sky130A

.subckt x3rd_3_OTA_flat vcc vss vo3 vd3 vd4 vb vd1
X0 a_1091_5624# vd4.t0 a_n515_844.t11 vss.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=17400,658 d=17400,658
X1 vcc.t15 a_n515_2006.t2 a_n515_2006.t3 vcc.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X2 vcc.t9 a_n515_844.t0 a_n515_844.t1 vcc.t8 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=29000,1116 d=14500,558
X3 a_1091_5624# vd4.t1 a_n515_844.t10 vss.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=34800,1316 d=17400,658
X4 a_n515_844.t9 vd4.t2 a_1091_5624# vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=34800,1316
X5 a_n515_2006.t7 a_n515_2006.t6 vcc.t14 vcc.t6 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=29000,1116
X6 a_n515_844.t7 a_n515_844.t6 vcc.t7 vcc.t6 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=29000,1116
X7 a_1091_5624# vd3.t0 a_n515_2006.t10 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=17400,658 d=17400,658
X8 vcc.t13 a_n515_2006.t4 a_n515_2006.t5 vcc.t8 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=29000,1116 d=14500,558
X9 a_3326_5370.t0 vo3.t0 vss.t4 sky130_fd_pr__res_xhigh_po_0p35 l=1.2
X10 vo3.t2 a_3898_4326# vss.t14 vss.t13 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X11 vss.t2 vb.t0 a_1091_5624# vss.t1 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=1.048143 ps=7.775429 w=5.5 l=1.5
**devattr s=63800,2316 d=31900,1158
X12 a_n515_844.t8 vd4.t3 a_1091_5624# vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=17400,658
X13 a_3898_4326# a_3898_4326# vss.t12 vss.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X14 vo3.t1 a_n515_844.t12 vcc.t5 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.6 l=0.35
**devattr s=30160,1156 d=30160,1156
X15 a_3326_5370.t1 vd1.t0 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X16 a_n515_844.t3 a_n515_844.t2 vcc.t3 vcc.t2 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X17 vcc.t1 a_n515_844.t4 a_n515_844.t5 vcc.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X18 a_1091_5624# vb.t1 vss.t9 vss.t1 sky130_fd_pr__nfet_01v8 ad=1.048143 pd=7.775429 as=0 ps=0 w=5.5 l=1.5
**devattr s=31900,1158 d=63800,2316
X19 a_1091_5624# vd3.t1 a_n515_2006.t0 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=34800,1316 d=17400,658
X20 a_n515_2006.t11 vd3.t2 a_1091_5624# vss.t15 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=17400,658
X21 a_n515_2006.t9 a_n515_2006.t8 vcc.t12 vcc.t2 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X22 a_n515_2006.t1 vd3.t3 a_1091_5624# vss.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=34800,1316
X23 a_3898_4326# a_n515_2006.t12 vcc.t11 vcc.t10 sky130_fd_pr__pfet_01v8_lvt ad=0.754 pd=5.78 as=0 ps=0 w=2.6 l=0.35
**devattr s=30160,1156 d=30160,1156
R0 vd4.n0 vd4.t2 82.3324
R1 vd4.n1 vd4.t3 81.6762
R2 vd4.n0 vd4.t0 81.6762
R3 vd4.n2 vd4.t1 81.4249
R4 vd4 vd4.n2 1.4105
R5 vd4.n1 vd4.n0 0.573
R6 vd4.n2 vd4.n1 0.238
R7 a_n515_844.n9 a_n515_844.t12 387.31
R8 a_n515_844.n8 a_n515_844.t7 96.3265
R9 a_n515_844.n6 a_n515_844.t1 96.3265
R10 a_n515_844.n3 a_n515_844.n10 84.9005
R11 a_n515_844.n5 a_n515_844.t10 35.0874
R12 a_n515_844.n5 a_n515_844.t9 34.5007
R13 a_n515_844.n9 a_n515_844.t6 32.649
R14 a_n515_844.t6 a_n515_844.n8 28.9361
R15 a_n515_844.n6 a_n515_844.n7 0.971171
R16 a_n515_844.n11 a_n515_844.n5 28.9205
R17 a_n515_844.n2 a_n515_844.t4 13.2766
R18 a_n515_844.t2 a_n515_844.n3 28.1453
R19 a_n515_844.t0 a_n515_844.n7 13.4238
R20 a_n515_844.n10 a_n515_844.t5 11.4265
R21 a_n515_844.n10 a_n515_844.t3 11.4265
R22 a_n515_844.n7 a_n515_844.n0 7.07514
R23 a_n515_844.n0 a_n515_844.n1 2.67922
R24 a_n515_844.t11 a_n515_844.n11 5.8005
R25 a_n515_844.n11 a_n515_844.t8 5.8005
R26 a_n515_844.n2 a_n515_844.n1 1.64285
R27 a_n515_844.n4 a_n515_844.n6 5.19734
R28 a_n515_844.n5 a_n515_844.n3 3.73846
R29 a_n515_844.n0 a_n515_844.n9 3.7305
R30 a_n515_844.n4 a_n515_844.n8 3.46037
R31 a_n515_844.n2 a_n515_844.n3 1.08359
R32 a_n515_844.n5 a_n515_844.n4 1.8052
R33 a_n515_844.t2 a_n515_844.n1 27.348
R34 vss.n28 vss.t7 102059
R35 vss.n77 vss.n12 12277.7
R36 vss.n77 vss.n13 12277.7
R37 vss.n85 vss.n12 12277.7
R38 vss.n85 vss.n13 12277.7
R39 vss.n28 vss.t6 11303
R40 vss.n74 vss.n9 6732.77
R41 vss.n87 vss.n9 6732.77
R42 vss.n74 vss.n10 6732.77
R43 vss.n87 vss.n10 6732.77
R44 vss.n31 vss.n19 4519.41
R45 vss.n49 vss.n19 4519.41
R46 vss.n31 vss.n20 4519.41
R47 vss.n49 vss.n20 4519.41
R48 vss.n39 vss.n25 3412.74
R49 vss.n37 vss.n25 3412.74
R50 vss.n39 vss.n26 3406.94
R51 vss.n37 vss.n26 3406.94
R52 vss.n32 vss.n28 3098.73
R53 vss.n46 vss.n21 1960.34
R54 vss.t6 vss.t10 1638.37
R55 vss.t7 vss.n11 1448.78
R56 vss.n27 vss.t15 847.806
R57 vss.t10 vss.n27 790.569
R58 vss.n78 vss.n15 588.515
R59 vss.n83 vss.n15 512.625
R60 vss.n76 vss.n50 462.808
R61 vss.n50 vss.n18 459.478
R62 vss.t3 vss.t8 381.233
R63 vss.n86 vss.n11 332.123
R64 vss.t0 vss.n85 301.05
R65 vss.n49 vss.n48 292.5
R66 vss.n50 vss.n49 292.5
R67 vss.n31 vss.n30 292.5
R68 vss.n32 vss.n31 292.5
R69 vss.n72 vss.n53 270.709
R70 vss.n76 vss.n75 257.209
R71 vss.n51 vss.t5 197.276
R72 vss.t15 vss.n11 189.595
R73 vss.t8 vss.t1 168.976
R74 vss.n38 vss.t13 149.831
R75 vss.n30 vss.n29 149.538
R76 vss.n38 vss.t11 146.5
R77 vss.t13 vss.n33 135.679
R78 vss.n29 vss.n21 126.4
R79 vss.n84 vss.n14 113.412
R80 vss.n84 vss.n83 109.558
R81 vss.n79 vss.n17 105.023
R82 vss.n35 vss.n26 97.5005
R83 vss.n26 vss.n18 97.5005
R84 vss.n34 vss.n25 97.5005
R85 vss.n33 vss.n25 97.5005
R86 vss.n23 vss.t14 89.2217
R87 vss.n23 vss.t12 89.0693
R88 vss.t4 vss.n18 80.7421
R89 vss.n36 vss.n34 73.0981
R90 vss.n37 vss.n36 65.0005
R91 vss.n38 vss.n37 65.0005
R92 vss.n40 vss.n39 65.0005
R93 vss.n39 vss.n38 65.0005
R94 vss.t11 vss.t4 57.4352
R95 vss.n36 vss.n35 56.241
R96 vss.n33 vss.n32 50.7761
R97 vss.n88 vss.n87 48.7505
R98 vss.n87 vss.n86 48.7505
R99 vss.n74 vss.n73 48.7505
R100 vss.n75 vss.n74 48.7505
R101 vss.t5 vss.n11 44.117
R102 vss.n75 vss.t3 38.2903
R103 vss.n41 vss.n20 34.4123
R104 vss.t4 vss.n20 34.4123
R105 vss.n29 vss.n19 34.4123
R106 vss.t4 vss.n19 34.4123
R107 vss.n14 vss.n8 34.0706
R108 vss.n55 vss.n10 32.5005
R109 vss.t1 vss.n10 32.5005
R110 vss.n59 vss.n9 32.5005
R111 vss.t1 vss.n9 32.5005
R112 vss.n45 vss.n22 30.4707
R113 vss.n59 vss.n58 28.0594
R114 vss.n71 vss.n70 24.7516
R115 vss.n54 vss.n8 24.4644
R116 vss.n30 vss.n24 20.517
R117 vss.n81 vss.n13 20.1729
R118 vss.n27 vss.n13 20.1729
R119 vss.n54 vss.n12 20.1729
R120 vss.n51 vss.n12 20.1729
R121 vss.n34 vss.n24 20.0772
R122 vss.n60 vss.n7 19.4026
R123 vss.n58 vss.n52 19.2005
R124 vss.n85 vss.n84 18.8715
R125 vss.n78 vss.n77 18.8715
R126 vss.n77 vss.n76 18.8715
R127 vss.n72 vss.n71 17.1218
R128 vss.n89 vss.n7 16.4046
R129 vss.n88 vss.n8 16.1396
R130 vss.t1 vss.n51 14.9835
R131 vss.n3 vss.n2 14.0913
R132 vss.n7 vss.n6 12.7191
R133 vss.n47 vss.n45 9.67855
R134 vss.n62 vss.n53 9.3005
R135 vss.n40 vss.n24 8.86924
R136 vss.n48 vss.n21 8.42977
R137 vss.n70 vss.n55 7.34725
R138 vss.n46 vss.n17 7.32557
R139 vss.n71 vss.n17 6.9983
R140 vss vss.n0 6.21349
R141 vss.n42 vss.n22 5.92892
R142 vss.n47 vss.n46 5.77749
R143 vss.n41 vss.n40 5.73359
R144 vss.n35 vss.n22 5.34506
R145 vss.n86 vss.t0 4.99482
R146 vss.n63 vss.n62 4.5005
R147 vss.n6 vss.n0 4.5005
R148 vss.n79 vss.n78 3.88247
R149 vss.n2 vss.t9 3.16414
R150 vss.n2 vss.t2 3.16414
R151 vss.n60 vss.n59 2.96471
R152 vss.n82 vss.n80 2.68449
R153 vss.n45 vss.n44 2.3255
R154 vss.n83 vss.n82 2.10165
R155 vss.n80 vss.n16 1.55874
R156 vss.n42 vss.n41 1.45132
R157 vss.n66 vss.n14 1.26099
R158 vss.n67 vss.n66 1.00227
R159 vss.n58 vss.n53 0.775237
R160 vss.n66 vss.n5 0.699787
R161 vss.n55 vss.n54 0.682157
R162 vss.n62 vss.n61 0.47062
R163 vss.n63 vss.n57 0.456098
R164 vss.n69 vss.n68 0.452003
R165 vss.n64 vss.n63 0.399937
R166 vss.n82 vss.n81 0.397733
R167 vss.n69 vss.n65 0.376108
R168 vss.n44 vss.n16 0.368932
R169 vss.n44 vss.n43 0.355
R170 vss.n61 vss.n4 0.350102
R171 vss.n57 vss.n1 0.344129
R172 vss.n68 vss.n67 0.326722
R173 vss.n65 vss.n64 0.311647
R174 vss.n80 vss.n79 0.3005
R175 vss.n62 vss.n56 0.272145
R176 vss.n48 vss.n47 0.250256
R177 vss.n93 vss.n92 0.227201
R178 vss.n73 vss.n72 0.224276
R179 vss.n56 vss.n52 0.221929
R180 vss.n68 vss.n5 0.221128
R181 vss.n91 vss.n4 0.220839
R182 vss.n67 vss.n3 0.216846
R183 vss.n90 vss.n5 0.209893
R184 vss.n81 vss.n15 0.180782
R185 vss.n90 vss.n89 0.133357
R186 vss.n70 vss.n69 0.126176
R187 vss.n43 vss.n42 0.122868
R188 vss.n43 vss.n23 0.118284
R189 vss.n61 vss.n60 0.107397
R190 vss.n92 vss.n91 0.0605
R191 vss vss.n93 0.048119
R192 vss.n61 vss.n57 0.0459545
R193 vss.n73 vss.n52 0.0452552
R194 vss.n1 vss.n0 0.0452485
R195 vss.n6 vss.n4 0.043226
R196 vss.n65 vss.n16 0.0382747
R197 vss.n89 vss.n88 0.027001
R198 vss.n64 vss.n56 0.0102403
R199 vss.n93 vss.n1 0.00456805
R200 vss.n92 vss.n3 0.00197929
R201 vss.n91 vss.n90 0.00155932
R202 a_n515_2006.n8 a_n515_2006.t12 387.724
R203 a_n515_2006.n4 a_n515_2006.t7 96.3265
R204 a_n515_2006.n7 a_n515_2006.t5 96.3265
R205 a_n515_2006.n0 a_n515_2006.n9 84.9005
R206 a_n515_2006.n3 a_n515_2006.t1 38.5285
R207 a_n515_2006.t0 a_n515_2006.n3 37.9091
R208 a_n515_2006.n3 a_n515_2006.t10 32.1034
R209 a_n515_2006.n5 a_n515_2006.n4 0.971171
R210 a_n515_2006.n7 a_n515_2006.n6 0.710684
R211 a_n515_2006.n0 a_n515_2006.t8 13.2778
R212 a_n515_2006.n1 a_n515_2006.n0 1.6868
R213 a_n515_2006.n6 a_n515_2006.t4 13.6521
R214 a_n515_2006.n5 a_n515_2006.t6 13.4238
R215 a_n515_2006.n1 a_n515_2006.t2 12.8838
R216 a_n515_2006.n9 a_n515_2006.t3 11.4265
R217 a_n515_2006.n9 a_n515_2006.t9 11.4265
R218 a_n515_2006.n0 a_n515_2006.n3 6.81377
R219 a_n515_2006.n3 a_n515_2006.n4 6.43072
R220 a_n515_2006.n2 a_n515_2006.n1 4.23945
R221 a_n515_2006.t10 a_n515_2006.t11 5.8005
R222 a_n515_2006.n8 a_n515_2006.n2 0.713738
R223 a_n515_2006.n2 a_n515_2006.n6 9.2977
R224 a_n515_2006.n5 a_n515_2006.n8 6.84764
R225 a_n515_2006.n7 a_n515_2006.n3 6.18407
R226 vcc.n60 vcc.n28 12420
R227 vcc.n60 vcc.n27 12420
R228 vcc.n58 vcc.n28 12416.5
R229 vcc.n58 vcc.n27 12416.5
R230 vcc.n64 vcc.n63 4698.77
R231 vcc.n16 vcc.n15 2071.76
R232 vcc.n23 vcc.n8 2071.76
R233 vcc.n20 vcc.n10 1443.53
R234 vcc.n20 vcc.n11 1443.53
R235 vcc.n47 vcc.n29 1037.16
R236 vcc.n16 vcc.n10 628.236
R237 vcc.n10 vcc.n8 628.236
R238 vcc.n13 vcc.n11 628.236
R239 vcc.n11 vcc.n9 628.236
R240 vcc.t0 vcc.t6 412.942
R241 vcc.t2 vcc.t8 412.942
R242 vcc.t6 vcc.n27 319.411
R243 vcc.t8 vcc.n28 315.507
R244 vcc.n47 vcc.n46 250.841
R245 vcc.n59 vcc.t2 208.423
R246 vcc.n59 vcc.t0 204.519
R247 vcc.n62 vcc.n61 177.656
R248 vcc.n21 vcc.t4 176.514
R249 vcc.t10 vcc.n21 176.514
R250 vcc.n15 vcc.n14 173.517
R251 vcc.n23 vcc.n22 173.517
R252 vcc.n62 vcc.n5 166.4
R253 vcc.n19 vcc.n18 153.976
R254 vcc.n19 vcc.n6 148.119
R255 vcc.n17 vcc.n12 124.802
R256 vcc.n39 vcc.t5 98.0045
R257 vcc.n39 vcc.t11 97.6911
R258 vcc.n24 vcc.n7 95.9841
R259 vcc.n63 vcc.n62 92.5809
R260 vcc.n36 vcc.n35 87.2408
R261 vcc.n42 vcc.n38 87.2408
R262 vcc.n32 vcc.n31 87.1446
R263 vcc.n52 vcc.n34 87.1446
R264 vcc.n48 vcc.n29 76.1836
R265 vcc.n18 vcc.n17 67.0123
R266 vcc.n18 vcc.n7 67.0123
R267 vcc.n12 vcc.n5 65.892
R268 vcc.n17 vcc.n16 61.6672
R269 vcc.n16 vcc.t4 61.6672
R270 vcc.n8 vcc.n7 61.6672
R271 vcc.t10 vcc.n8 61.6672
R272 vcc.n13 vcc.n5 61.6672
R273 vcc.n9 vcc.n6 61.6672
R274 vcc.n65 vcc.n4 57.3115
R275 vcc.n14 vcc.n13 54.8697
R276 vcc.n22 vcc.n9 54.8697
R277 vcc.n62 vcc.n25 41.9251
R278 vcc.n57 vcc.n2 35.1478
R279 vcc.n55 vcc.n29 34.0937
R280 vcc.n65 vcc.n64 24.2792
R281 vcc.n20 vcc.n19 18.5005
R282 vcc.n21 vcc.n20 18.5005
R283 vcc.n15 vcc.n12 18.5005
R284 vcc.n24 vcc.n23 18.5005
R285 vcc.n25 vcc.n24 18.273
R286 vcc.n61 vcc.n26 11.6663
R287 vcc.n31 vcc.t7 11.4265
R288 vcc.n31 vcc.t15 11.4265
R289 vcc.n34 vcc.t12 11.4265
R290 vcc.n34 vcc.t9 11.4265
R291 vcc.n35 vcc.t3 11.4265
R292 vcc.n35 vcc.t13 11.4265
R293 vcc.n38 vcc.t14 11.4265
R294 vcc.n38 vcc.t1 11.4265
R295 vcc.n37 vcc.n26 9.3005
R296 vcc.n68 vcc.n2 9.3005
R297 vcc.n55 vcc.n54 9.3005
R298 vcc.n49 vcc.n47 8.86797
R299 vcc.n62 vcc.n6 8.01848
R300 vcc.n70 vcc.n1 6.3755
R301 vcc.n48 vcc.n28 5.60656
R302 vcc.n27 vcc.n4 5.60656
R303 vcc.n14 vcc.t4 5.16575
R304 vcc.n22 vcc.t10 5.16575
R305 vcc.n43 vcc.n37 4.5005
R306 vcc.n54 vcc.n53 4.5005
R307 vcc.n69 vcc.n68 4.5005
R308 vcc.n45 vcc.n30 3.83011
R309 vcc.n63 vcc.n4 3.30373
R310 vcc.n40 vcc.n37 3.09113
R311 vcc.n61 vcc.n60 2.68166
R312 vcc.n60 vcc.n59 2.68166
R313 vcc.n58 vcc.n57 2.68166
R314 vcc.n59 vcc.n58 2.68166
R315 vcc.n51 vcc.n36 2.57239
R316 vcc.n68 vcc.n67 1.97251
R317 vcc.n54 vcc.n30 1.78308
R318 vcc.n42 vcc.n41 1.688
R319 vcc.n52 vcc.n51 1.60959
R320 vcc.n46 vcc.n26 1.45873
R321 vcc vcc.n70 1.43376
R322 vcc.n43 vcc.n42 1.27935
R323 vcc.n56 vcc.n55 1.19015
R324 vcc.n64 vcc.n2 1.05462
R325 vcc.n67 vcc.n66 1.039
R326 vcc.n44 vcc.n36 0.963107
R327 vcc.n67 vcc.n65 0.845955
R328 vcc.n68 vcc.n3 0.780009
R329 vcc.n40 vcc.n25 0.58175
R330 vcc.n32 vcc.n1 0.39076
R331 vcc.n33 vcc.n32 0.347903
R332 vcc.n53 vcc.n52 0.314461
R333 vcc.n57 vcc.n56 0.2565
R334 vcc.n41 vcc.n40 0.2505
R335 vcc.n50 vcc.n49 0.1505
R336 vcc.n46 vcc.n45 0.148119
R337 vcc.n69 vcc.n0 0.144487
R338 vcc.n41 vcc.n39 0.133423
R339 vcc.n49 vcc.n48 0.0776084
R340 vcc.n51 vcc.n50 0.0666765
R341 vcc.n45 vcc.n44 0.0638803
R342 vcc.n56 vcc.n3 0.0274565
R343 vcc.n54 vcc.n3 0.0266936
R344 vcc.n53 vcc.n33 0.0261494
R345 vcc vcc.n0 0.0216864
R346 vcc.n45 vcc.n37 0.0211422
R347 vcc.n44 vcc.n43 0.0197308
R348 vcc.n66 vcc.n1 0.0170584
R349 vcc.n50 vcc.n30 0.014395
R350 vcc.n33 vcc.n3 0.0121883
R351 vcc.n70 vcc.n69 0.00841139
R352 vcc.n66 vcc.n0 0.00129114
R353 vd3.n0 vd3.t3 81.6812
R354 vd3.n1 vd3.t2 81.6574
R355 vd3.n0 vd3.t0 81.6574
R356 vd3.n2 vd3.t1 81.4437
R357 vd3 vd3.n2 1.0755
R358 vd3.n2 vd3.n1 0.908
R359 vd3.n1 vd3.n0 0.573
R360 a_3326_5370.t0 a_3326_5370.t1 50.1091
R361 vo3.n0 vo3.t1 98.5661
R362 vo3.n0 vo3.t2 88.8259
R363 vo3.n1 vo3.t0 46.6411
R364 vo3.n1 vo3.n0 0.509181
R365 vo3 vo3.n1 0.267861
R366 vb.n0 vb.t1 69.2431
R367 vb.n0 vb.t0 68.768
R368 vb vb.n0 40.2939
R369 vd1 vd1.t0 0.121075
C0 vcc vo3 0.586239f
C1 a_3898_4326# vcc 0.836592f
C2 vd3 vcc 0.03196f
C3 vcc a_1091_5624# 0.101608f
C4 vd3 vb 0.10442f
C5 a_1091_5624# vb 0.545685f
C6 vd1 vo3 0.023381f
C7 vd4 a_3898_4326# 1.15e-20
C8 vd4 vd3 2.98724f
C9 a_3898_4326# vd1 0.002363f
C10 vcc vb 2.02e-19
C11 vd4 a_1091_5624# 1.05152f
C12 a_1091_5624# vd1 0.006984f
C13 a_3898_4326# vo3 0.159329f
C14 vd4 vcc 0.055614f
C15 vd3 a_3898_4326# 4.42e-20
C16 a_1091_5624# vo3 0.004168f
C17 a_3898_4326# a_1091_5624# 0.016974f
C18 vd4 vb 0.028439f
C19 vd3 a_1091_5624# 1.06971f
C20 vb vd1 0.036045f
C21 vd1 vss 9.14385f
C22 vd4 vss 5.653077f
C23 vd3 vss 5.6615f
C24 vo3 vss 2.14738f
C25 vb vss 4.13375f
C26 vcc vss 50.4443f
C27 a_3898_4326# vss 1.47495f
C28 a_1091_5624# vss 5.74998f
C29 vd1.t0 vss 25.0601f
C30 a_3326_5370.t1 vss 26.271801f
C31 a_3326_5370.t0 vss 0.028206f
C32 vd3.t3 vss 0.471581f
C33 vd3.t0 vss 0.471443f
C34 vd3.n0 vss 0.4652f
C35 vd3.t2 vss 0.471443f
C36 vd3.n1 vss 0.270746f
C37 vd3.t1 vss 0.470875f
C38 vd3.n2 vss 0.302202f
C39 vcc.n0 vss 0.035285f
C40 vcc.n1 vss 0.222321f
C41 vcc.n2 vss 0.941429f
C42 vcc.n3 vss 0.422066f
C43 vcc.n4 vss 0.052416f
C44 vcc.n5 vss 0.165753f
C45 vcc.n6 vss 0.054389f
C46 vcc.n7 vss 0.019349f
C47 vcc.n8 vss 0.012354f
C48 vcc.n9 vss 0.012354f
C49 vcc.t4 vss 0.169018f
C50 vcc.n10 vss 0.011983f
C51 vcc.n11 vss 0.011983f
C52 vcc.n12 vss 0.047323f
C53 vcc.n13 vss 0.012354f
C54 vcc.n15 vss 0.13217f
C55 vcc.n16 vss 0.012354f
C56 vcc.n17 vss 0.016164f
C57 vcc.n18 vss 0.011983f
C58 vcc.n19 vss 0.012621f
C59 vcc.n20 vss 0.012814f
C60 vcc.n21 vss 0.157127f
C61 vcc.t10 vss 0.169018f
C62 vcc.n23 vss 0.13217f
C63 vcc.n24 vss 0.059919f
C64 vcc.n25 vss 0.041263f
C65 vcc.n26 vss 0.011792f
C66 vcc.n27 vss 1.1135f
C67 vcc.n28 vss 1.13751f
C68 vcc.t6 vss 2.10593f
C69 vcc.t0 vss 1.77403f
C70 vcc.n29 vss 1.1934f
C71 vcc.n30 vss 0.43099f
C72 vcc.t7 vss 0.00668f
C73 vcc.t15 vss 0.00668f
C74 vcc.n31 vss 0.014478f
C75 vcc.n32 vss 0.45615f
C76 vcc.n33 vss 0.203805f
C77 vcc.t12 vss 0.00668f
C78 vcc.t9 vss 0.00668f
C79 vcc.n34 vss 0.014478f
C80 vcc.t3 vss 0.00668f
C81 vcc.t13 vss 0.00668f
C82 vcc.n35 vss 0.014537f
C83 vcc.n36 vss 0.236013f
C84 vcc.n37 vss 0.139136f
C85 vcc.t14 vss 0.00668f
C86 vcc.t1 vss 0.00668f
C87 vcc.n38 vss 0.014537f
C88 vcc.t5 vss 0.026632f
C89 vcc.t11 vss 0.026418f
C90 vcc.n39 vss 0.13963f
C91 vcc.n40 vss 0.219712f
C92 vcc.n41 vss 0.046033f
C93 vcc.n42 vss 0.204361f
C94 vcc.n43 vss 0.065493f
C95 vcc.n44 vss 0.049537f
C96 vcc.n45 vss 0.169314f
C97 vcc.n46 vss 0.232881f
C98 vcc.n47 vss 0.277736f
C99 vcc.n48 vss 0.075638f
C100 vcc.n49 vss 0.008872f
C101 vcc.n50 vss 0.055054f
C102 vcc.n51 vss 0.281487f
C103 vcc.n52 vss 0.702843f
C104 vcc.n53 vss 0.185534f
C105 vcc.n54 vss 0.70362f
C106 vcc.n55 vss 0.91754f
C107 vcc.n56 vss 0.037595f
C108 vcc.n57 vss 0.920673f
C109 vcc.n58 vss 0.110557f
C110 vcc.t8 vss 2.09537f
C111 vcc.t2 vss 1.78524f
C112 vcc.n59 vss 1.18642f
C113 vcc.n60 vss 0.110589f
C114 vcc.n61 vss 0.170722f
C115 vcc.n62 vss 0.376561f
C116 vcc.n63 vss 0.090974f
C117 vcc.n64 vss 0.111214f
C118 vcc.n65 vss 0.070554f
C119 vcc.n66 vss 0.070038f
C120 vcc.n67 vss 0.120865f
C121 vcc.n68 vss 0.45792f
C122 vcc.n69 vss 0.013976f
C123 vcc.n70 vss 0.001968f
C124 a_n515_2006.n0 vss 1.46343f
C125 a_n515_2006.n1 vss 0.936679f
C126 a_n515_2006.n2 vss 1.29294f
C127 a_n515_2006.n3 vss 5.4296f
C128 a_n515_2006.n4 vss 0.906852f
C129 a_n515_2006.n5 vss 0.620305f
C130 a_n515_2006.n6 vss 0.742801f
C131 a_n515_2006.n7 vss 0.763129f
C132 a_n515_2006.n8 vss 1.26286f
C133 a_n515_2006.t1 vss 0.150208f
C134 a_n515_2006.t7 vss 0.080806f
C135 a_n515_2006.t12 vss 0.127287f
C136 a_n515_2006.t4 vss 1.5052f
C137 a_n515_2006.t5 vss 0.080806f
C138 a_n515_2006.t8 vss 1.48973f
C139 a_n515_2006.t3 vss 0.021976f
C140 a_n515_2006.t9 vss 0.021976f
C141 a_n515_2006.n9 vss 0.044771f
C142 a_n515_2006.t2 vss 1.48363f
C143 a_n515_2006.t6 vss 1.49909f
C144 a_n515_2006.t10 vss 0.109556f
C145 a_n515_2006.t11 vss 0.026371f
C146 a_n515_2006.t0 vss 0.139993f
C147 a_n515_844.n0 vss 1.17962f
C148 a_n515_844.n1 vss 1.22804f
C149 a_n515_844.n2 vss 0.281253f
C150 a_n515_844.n3 vss 1.29217f
C151 a_n515_844.n4 vss 1.58696f
C152 a_n515_844.n5 vss 3.86796f
C153 a_n515_844.n6 vss 1.02899f
C154 a_n515_844.n7 vss 0.64178f
C155 a_n515_844.t8 vss 0.026714f
C156 a_n515_844.t7 vss 0.081856f
C157 a_n515_844.n8 vss 0.711803f
C158 a_n515_844.t12 vss 0.12612f
C159 a_n515_844.t6 vss 1.63702f
C160 a_n515_844.n9 vss 1.63593f
C161 a_n515_844.t5 vss 0.022262f
C162 a_n515_844.t3 vss 0.022262f
C163 a_n515_844.n10 vss 0.045353f
C164 a_n515_844.t4 vss 1.50909f
C165 a_n515_844.t2 vss 1.52061f
C166 a_n515_844.t0 vss 1.51857f
C167 a_n515_844.t1 vss 0.081856f
C168 a_n515_844.t10 vss 0.129668f
C169 a_n515_844.t9 vss 0.118903f
C170 a_n515_844.n11 vss 0.078484f
C171 a_n515_844.t11 vss 0.026714f
C172 vd4.t2 vss 0.471605f
C173 vd4.t0 vss 0.473171f
C174 vd4.n0 vss 0.511022f
C175 vd4.t3 vss 0.473171f
C176 vd4.n1 vss 0.249669f
C177 vd4.t1 vss 0.469223f
C178 vd4.n2 vss 0.251842f
.ends

