** sch_path: /home/zerotoasic/Project_tinytape/xschem/Projects/tinytape/OTA/OTA_tinytape/layout
*+ schs/BGR_BJT_stage2.sch
.subckt BGR_BJT_stage2 vb vcc vss vref0 vr vb1
*.PININFO vb:O vcc:I vss:I vref0:I vr:I vb1:O
XM4 net1 net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM5 net2 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM6 vb1 net3 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM7 net3 net3 vb1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM10 net2 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM11 net3 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM12 vb vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM16 net4 net5 vb1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM15 net5 net5 net4 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM14 net5 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM19 vb net6 net4 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM18 net6 net6 vb vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM17 net6 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM1 net2 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM2 net2 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM3 net2 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM8 net3 net3 vb1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM9 net3 net3 vb1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM13 net3 net3 vb1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM20 net5 net5 net4 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM21 net5 net5 net4 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM22 net5 net5 net4 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM23 net6 net6 vb vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM24 net6 net6 vb vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM25 net6 net6 vb vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
.ends
.end
