* NGSPICE file created from 3_OTA_flat.ext - technology: sky130A

.subckt x3_OTA_flat vo3 vin_p vin_n vcc vss
X0 a_9040_n3397# 2nd_3_OTA_0.vd3.t12 a_7434_495.t3 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=34800,1316 d=17400,658
X1 a_n1236_n9479.t47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X2 a_7434_1657.t11 2nd_3_OTA_0.vd4.t8 a_9040_n3397# vss.t51 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=17400,658
X3 2nd_3_OTA_0.vd3.t2 2nd_3_OTA_0.vd2.t5 a_n1050_166.t10 vcc.t27 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X4 2nd_3_OTA_0.vd2.t0 vin_p.t0 a_n10077_1624# vss.t11 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X5 vo3.t0 a_7434_1657.t12 vcc.t14 vcc.t13 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.6 l=0.35
**devattr s=30160,1156 d=30160,1156
X6 a_n1236_n9479.t46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X7 a_n1236_n9479.t45 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 OTA_vref_0.OTA_vref_stage2_0.vref0.t32 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X8 a_7434_1657.t1 a_7434_1657.t0 vcc.t12 vcc.t11 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X9 a_7434_495.t5 a_7434_495.t4 vcc.t49 vcc.t9 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=29000,1116
X10 2nd_3_OTA_0.vb1.t5 a_2382_n6868# a_2470_n7958# vss.t22 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X11 a_n1236_n9479.t44 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X12 a_2382_n8158# OTA_vref_0.OTA_vref_stage2_0.vr.t20 vcc.t36 vcc.t35 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X13 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 a_n1236_n9479.t43 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X14 a_11847_n1701# a_11847_n1701# vss.t29 vss.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X15 vss.t62 2nd_3_OTA_0.vd3.t4 2nd_3_OTA_0.vd3.t5 vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X16 a_11275_n2439.t1 3rd_3_OTA_0.vd1 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X17 2nd_3_OTA_0.vd2.t2 2nd_3_OTA_0.vd2.t1 vcc.t43 vcc.t41 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X18 vss.t7 a_n1236_n9479.t30 a_n1236_n9479.t31 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X19 OTA_vref_0.vb a_2382_n4288# a_2382_n4288# vss.t50 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X20 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 a_n1236_n9479.t42 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X21 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 a_n1236_n9479.t41 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X22 vss.t6 vss.t30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X23 2nd_3_OTA_0.vd1.t1 2nd_3_OTA_0.vd2.t1 vcc.t42 vcc.t41 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X24 a_n10077_1624# vin_p.t1 2nd_3_OTA_0.vd2.t4 vss.t64 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X25 a_7434_1657.t5 a_7434_1657.t4 vcc.t10 vcc.t9 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=29000,1116
X26 vss.t39 a_n1236_n9479.t28 a_n1236_n9479.t29 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X27 a_11847_n1701# a_7434_495.t12 vcc.t48 vcc.t47 sky130_fd_pr__pfet_01v8_lvt ad=0.754 pd=5.78 as=0 ps=0 w=2.6 l=0.35
**devattr s=30160,1156 d=30160,1156
X28 a_7434_495.t2 2nd_3_OTA_0.vd3.t13 a_9040_n3397# vss.t51 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=17400,658
X29 a_2382_n6868# a_2382_n6868# 2nd_3_OTA_0.vb1.t4 vss.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X30 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 a_n1236_n9479.t40 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X31 OTA_vref_0.OTA_vref_stage2_0.vr.t19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X32 2nd_3_OTA_0.vd3.t9 2nd_3_OTA_0.vd3.t8 vss.t61 vss.t56 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X33 vcc.t8 a_7434_1657.t2 a_7434_1657.t3 vcc.t7 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X34 a_2470_n7958# a_2382_n8158# a_2382_n8158# vss.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X35 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 a_n1236_n9479.t39 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X36 OTA_vref_0.OTA_vref_stage2_0.vr.t18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X37 a_n1050_166.t9 2nd_3_OTA_0.vd2.t6 2nd_3_OTA_0.vd3.t3 vcc.t30 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X38 a_2382_n6868# a_2382_n6868# 2nd_3_OTA_0.vb1.t3 vss.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X39 vcc.t6 a_7434_1657.t6 a_7434_1657.t7 vcc.t5 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=29000,1116 d=14500,558
X40 a_2382_n4288# a_2382_n4288# OTA_vref_0.vb vss.t49 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=5800,258 d=5800,258
X41 a_n1236_n9479.t38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X42 a_n1050_166.t0 2nd_3_OTA_0.vb1.t6 vcc.t1 vcc.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=81200,2916
X43 2nd_3_OTA_0.vd4.t9 3rd_3_OTA_0.vd1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X44 vss.t25 a_n1236_n9479.t26 a_n1236_n9479.t27 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X45 OTA_vref_0.OTA_vref_stage2_0.vr.t17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X46 OTA_vref_0.OTA_vref_stage2_0.vr.t16 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X47 OTA_vref_0.OTA_vref_stage2_0.vr.t3 OTA_vref_0.OTA_vref_stage2_0.vr.t2 vcc.t33 vcc.t32 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=2900,158 d=5800,316
X48 vss.t60 2nd_3_OTA_0.vd3.t14 2nd_3_OTA_0.vd4.t6 vss.t54 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X49 2nd_3_OTA_0.vb1.t2 a_2382_n6868# a_2382_n6868# vss.t19 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X50 vcc.t26 2nd_3_OTA_0.vb1.t7 a_n1050_166.t3 vcc.t25 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X51 vss.t38 a_n1236_n9479.t24 a_n1236_n9479.t25 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X52 a_9040_n3397# 2nd_3_OTA_0.vd4.t10 a_7434_1657.t10 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=34800,1316 d=17400,658
X53 OTA_vref_0.vb a_2382_n4288# a_2470_n5378# vss.t48 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X54 a_2382_n5578# OTA_vref_0.OTA_vref_stage2_0.vr.t21 vcc.t22 vcc.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X55 vss.t23 a_n1236_n9479.t22 a_n1236_n9479.t23 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X56 vss.t40 a_n1236_n9479.t20 a_n1236_n9479.t21 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X57 a_n1050_166.t6 2nd_3_OTA_0.vd1.t4 2nd_3_OTA_0.vd4.t2 vcc.t30 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X58 vss.t17 a_n1236_n9479.t18 a_n1236_n9479.t19 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X59 a_n10077_1624# vin_n.t0 2nd_3_OTA_0.vd1.t2 vss.t65 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X60 a_2470_n7958# a_2382_n8158# OTA_vref_0.OTA_vref_stage2_0.vref0.t0 vss.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X61 vcc.t3 2nd_3_OTA_0.vb1.t8 a_n1050_166.t1 vcc.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=81200,2916 d=40600,1458
X62 a_n1050_166.t11 2nd_3_OTA_0.vd1.t5 2nd_3_OTA_0.vd4.t7 vcc.t40 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X63 2nd_3_OTA_0.vd3.t7 2nd_3_OTA_0.vd3.t6 vss.t59 vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X64 a_n1236_n9479.t17 a_n1236_n9479.t16 vss.t32 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X65 a_2382_n4288# a_2382_n4288# OTA_vref_0.vb vss.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=5800,258 d=5800,258
X66 OTA_vref_0.OTA_vref_stage2_0.vr.t15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X67 vss.t31 a_n1236_n9479.t14 a_n1236_n9479.t15 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X68 a_n1050_166.t8 2nd_3_OTA_0.vd2.t7 2nd_3_OTA_0.vd3.t1 vcc.t40 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X69 a_n1236_n9479.t13 a_n1236_n9479.t12 vss.t44 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X70 a_2470_n5378# a_2382_n5578# a_2382_n5578# vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X71 vcc.t24 OTA_vref_0.OTA_vref_stage2_0.vr.t22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 vcc.t23 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X72 vss.t58 2nd_3_OTA_0.vd3.t15 2nd_3_OTA_0.vd4.t5 vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X73 OTA_vref_0.OTA_vref_stage2_0.vr.t14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X74 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 OTA_vref_0.OTA_vref_stage2_0.vr.t13 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X75 OTA_vref_0.OTA_vref_stage2_0.vr.t12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X76 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 OTA_vref_0.OTA_vref_stage2_0.vr.t11 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X77 a_7434_1657.t9 2nd_3_OTA_0.vd4.t11 a_9040_n3397# vss.t41 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=34800,1316
X78 2nd_3_OTA_0.vd3.t0 2nd_3_OTA_0.vd2.t8 a_n1050_166.t7 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X79 a_2382_n8158# a_2382_n8158# a_2470_n7958# vss.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X80 2nd_3_OTA_0.vd1.t3 vin_n.t1 a_n10077_1624# vss.t66 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X81 a_2382_n5578# a_2382_n5578# a_2470_n5378# vss.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X82 a_7434_495.t11 a_7434_495.t10 vcc.t46 vcc.t11 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X83 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 a_n1236_n9479.t37 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X84 OTA_vref_0.vb a_2382_n4288# a_2382_n4288# vss.t46 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=11600,516
X85 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 OTA_vref_0.OTA_vref_stage2_0.vr.t10 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X86 a_n1050_166.t5 2nd_3_OTA_0.vb1.t9 vcc.t29 vcc.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 OTA_vref_0.OTA_vref_stage2_0.vr.t23 vcc.t20 vcc.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=11600,516
X88 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 OTA_vref_0.OTA_vref_stage2_0.vr.t9 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X89 a_2470_n5378# a_2382_n5578# 2nd_3_OTA_0.vb1.t0 vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X90 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 OTA_vref_0.OTA_vref_stage2_0.vr.t8 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X91 a_2382_n6868# OTA_vref_0.OTA_vref_stage2_0.vr.t24 vcc.t18 vcc.t17 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X92 a_n1236_n9479.t11 a_n1236_n9479.t10 vss.t45 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X93 a_2470_n7958# a_2382_n8158# a_2382_n8158# vss.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X94 vcc.t45 a_7434_495.t6 a_7434_495.t7 vcc.t7 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X95 2nd_3_OTA_0.vd4.t4 2nd_3_OTA_0.vd3.t16 vss.t57 vss.t56 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X96 a_n1236_n9479.t9 a_n1236_n9479.t8 vss.t42 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X97 a_n1236_n9479.t7 a_n1236_n9479.t6 vss.t8 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X98 vo3.t2 a_11847_n1701# vss.t27 vss.t26 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X99 a_9040_n3397# 2nd_3_OTA_0.vd4.t12 a_7434_1657.t8 vss.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=17400,658 d=17400,658
X100 vss.t55 2nd_3_OTA_0.vd3.t10 2nd_3_OTA_0.vd3.t11 vss.t54 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X101 a_2382_n8158# a_2382_n8158# a_2470_n7958# vss.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X102 a_n1236_n9479.t5 a_n1236_n9479.t4 vss.t63 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X103 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 OTA_vref_0.OTA_vref_stage2_0.vr.t7 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X104 vcc.t39 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd1.t0 vcc.t37 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X105 vcc.t34 OTA_vref_0.OTA_vref_stage2_0.vr.t0 OTA_vref_0.OTA_vref_stage2_0.vr.t1 vcc.t32 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=5800,316 d=2900,158
X106 a_n1236_n9479.t36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X107 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 a_n1236_n9479.t35 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X108 a_2382_n5578# a_2382_n5578# a_2470_n5378# vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X109 a_n1236_n9479.t3 a_n1236_n9479.t2 vss.t43 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X110 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 a_n1236_n9479.t34 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X111 2nd_3_OTA_0.vd4.t0 2nd_3_OTA_0.vd1.t6 a_n1050_166.t2 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X112 2nd_3_OTA_0.vb1.t1 a_2382_n6868# a_2382_n6868# vss.t18 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X113 OTA_vref_0.vb OTA_vref_0.OTA_vref_stage2_0.vr.t25 vcc.t31 vcc.t15 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X114 2nd_3_OTA_0.vd4.t1 2nd_3_OTA_0.vd1.t7 a_n1050_166.t4 vcc.t27 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X115 vcc.t38 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd2.t3 vcc.t37 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X116 vcc.t44 a_7434_495.t8 a_7434_495.t9 vcc.t5 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=29000,1116 d=14500,558
X117 a_9040_n3397# OTA_vref_0.vb vss.t37 vss.t33 sky130_fd_pr__nfet_01v8 ad=1.048143 pd=7.775429 as=0 ps=0 w=5.5 l=1.5
**devattr s=31900,1158 d=63800,2316
X118 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 OTA_vref_0.OTA_vref_stage2_0.vr.t6 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X119 2nd_3_OTA_0.vd4.t3 2nd_3_OTA_0.vd3.t17 vss.t53 vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X120 a_n1236_n9479.t33 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X121 a_n10077_1624# OTA_vref_0.vb vss.t36 vss.t35 sky130_fd_pr__nfet_01v8 ad=0.483333 pd=3.526667 as=0 ps=0 w=3 l=5
**devattr s=34800,1316 d=34800,1316
X122 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 OTA_vref_0.OTA_vref_stage2_0.vr.t5 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X123 a_9040_n3397# 2nd_3_OTA_0.vd3.t18 a_7434_495.t1 vss.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=17400,658 d=17400,658
X124 a_n1236_n9479.t32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X125 a_11275_n2439.t0 vo3.t1 vss.t24 sky130_fd_pr__res_xhigh_po_0p35 l=1.2
X126 a_2382_n4288# OTA_vref_0.OTA_vref_stage2_0.vr.t26 vcc.t16 vcc.t15 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X127 OTA_vref_0.OTA_vref_stage2_0.vr.t4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X128 a_7434_495.t0 2nd_3_OTA_0.vd3.t19 a_9040_n3397# vss.t41 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=34800,1316
X129 vss.t34 OTA_vref_0.vb a_9040_n3397# vss.t33 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=1.048143 ps=7.775429 w=5.5 l=1.5
**devattr s=63800,2316 d=31900,1158
X130 a_2470_n5378# a_2382_n5578# a_2382_n5578# vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X131 a_n1236_n9479.t1 a_n1236_n9479.t0 vss.t67 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
R0 2nd_3_OTA_0.vd3.n0 2nd_3_OTA_0.vd3.t19 81.6812
R1 2nd_3_OTA_0.vd3.n0 2nd_3_OTA_0.vd3.t13 81.6574
R2 2nd_3_OTA_0.vd3.n0 2nd_3_OTA_0.vd3.t18 81.6574
R3 2nd_3_OTA_0.vd3 2nd_3_OTA_0.vd3.t12 81.4437
R4 2nd_3_OTA_0.vd3.n2 2nd_3_OTA_0.vd3.t9 60.3532
R5 2nd_3_OTA_0.vd3.n1 2nd_3_OTA_0.vd3.t11 60.3532
R6 2nd_3_OTA_0.vd3.n3 2nd_3_OTA_0.vd3.n10 48.5755
R7 2nd_3_OTA_0.vd3.n5 2nd_3_OTA_0.vd3.t1 19.1315
R8 2nd_3_OTA_0.vd3.n5 2nd_3_OTA_0.vd3.t2 18.308
R9 2nd_3_OTA_0.vd3.n5 2nd_3_OTA_0.vd3.n6 16.2724
R10 2nd_3_OTA_0.vd3.n13 2nd_3_OTA_0.vd3.n1 14.6534
R11 2nd_3_OTA_0.vd3.n10 2nd_3_OTA_0.vd3.t5 11.6005
R12 2nd_3_OTA_0.vd3.n10 2nd_3_OTA_0.vd3.t7 11.6005
R13 2nd_3_OTA_0.vd3 2nd_3_OTA_0.vd3.n1 11.2227
R14 2nd_3_OTA_0.vd3.n3 2nd_3_OTA_0.vd3.n7 8.08817
R15 2nd_3_OTA_0.vd3 2nd_3_OTA_0.vd3.n2 7.9105
R16 2nd_3_OTA_0.vd3.n8 2nd_3_OTA_0.vd3.t8 3.58326
R17 2nd_3_OTA_0.vd3.n9 2nd_3_OTA_0.vd3.t15 3.58326
R18 2nd_3_OTA_0.vd3.n11 2nd_3_OTA_0.vd3.t17 3.58326
R19 2nd_3_OTA_0.vd3.n12 2nd_3_OTA_0.vd3.t10 3.58326
R20 2nd_3_OTA_0.vd3.n8 2nd_3_OTA_0.vd3.t16 3.58267
R21 2nd_3_OTA_0.vd3.n9 2nd_3_OTA_0.vd3.t4 3.58267
R22 2nd_3_OTA_0.vd3.n11 2nd_3_OTA_0.vd3.t6 3.58267
R23 2nd_3_OTA_0.vd3.n12 2nd_3_OTA_0.vd3.t14 3.58267
R24 2nd_3_OTA_0.vd3.n4 2nd_3_OTA_0.vd3.n13 3.54985
R25 2nd_3_OTA_0.vd3.n7 2nd_3_OTA_0.vd3.n5 2.67636
R26 2nd_3_OTA_0.vd3.n1 2nd_3_OTA_0.vd3.n12 2.60735
R27 2nd_3_OTA_0.vd3.n2 2nd_3_OTA_0.vd3.n8 2.58162
R28 2nd_3_OTA_0.vd3 2nd_3_OTA_0.vd3.n0 2.5555
R29 2nd_3_OTA_0.vd3 2nd_3_OTA_0.vd3.n7 2.29713
R30 2nd_3_OTA_0.vd3.n6 2nd_3_OTA_0.vd3.t3 1.90483
R31 2nd_3_OTA_0.vd3.n6 2nd_3_OTA_0.vd3.t0 1.90483
R32 2nd_3_OTA_0.vd3.n2 2nd_3_OTA_0.vd3.n4 1.69798
R33 2nd_3_OTA_0.vd3.n13 2nd_3_OTA_0.vd3.n11 1.61224
R34 2nd_3_OTA_0.vd3.n4 2nd_3_OTA_0.vd3.n9 1.61224
R35 2nd_3_OTA_0.vd3.n4 2nd_3_OTA_0.vd3.n3 1.22519
R36 a_7434_495.n8 a_7434_495.t12 387.724
R37 a_7434_495.n7 a_7434_495.t9 96.3265
R38 a_7434_495.n4 a_7434_495.t5 96.3265
R39 a_7434_495.n0 a_7434_495.n9 84.9005
R40 a_7434_495.n3 a_7434_495.t0 38.5275
R41 a_7434_495.t3 a_7434_495.n3 37.908
R42 a_7434_495.n3 a_7434_495.n10 32.1023
R43 a_7434_495.n4 a_7434_495.n5 0.971171
R44 a_7434_495.n7 a_7434_495.n6 0.710684
R45 a_7434_495.n0 a_7434_495.t10 13.2778
R46 a_7434_495.n1 a_7434_495.n0 1.6868
R47 a_7434_495.n6 a_7434_495.t8 13.6521
R48 a_7434_495.n1 a_7434_495.t6 12.8838
R49 a_7434_495.t4 a_7434_495.n5 13.4238
R50 a_7434_495.n9 a_7434_495.t7 11.4265
R51 a_7434_495.n9 a_7434_495.t11 11.4265
R52 a_7434_495.n0 a_7434_495.n3 6.81377
R53 a_7434_495.n3 a_7434_495.n4 6.43072
R54 a_7434_495.n2 a_7434_495.n1 4.23945
R55 a_7434_495.n10 a_7434_495.t1 5.8005
R56 a_7434_495.n10 a_7434_495.t2 5.8005
R57 a_7434_495.n8 a_7434_495.n2 0.713738
R58 a_7434_495.n2 a_7434_495.n6 9.2977
R59 a_7434_495.n5 a_7434_495.n8 6.84764
R60 a_7434_495.n7 a_7434_495.n3 6.18407
R61 vss.n53 vss.t52 6.51798e+06
R62 vss.n311 vss.n57 5.4843e+06
R63 vss.n57 vss.n54 3.3e+06
R64 vss.n54 vss.n53 2.376e+06
R65 vss.n313 vss.n312 1.23016e+06
R66 vss.n313 vss.n54 402600
R67 vss.n312 vss.n311 354428
R68 vss.n367 vss.n315 156933
R69 vss.n465 vss.n6 147329
R70 vss.n336 vss.n315 114006
R71 vss.n466 vss.n465 72897.2
R72 vss.t52 vss.n6 36497.6
R73 vss.n467 vss.n466 31912.6
R74 vss.n463 vss.n7 27614.8
R75 vss.n463 vss.n8 27609
R76 vss.n450 vss.n7 27609
R77 vss.n450 vss.n8 27603.2
R78 vss.n443 vss.n33 26954.2
R79 vss.n422 vss.n33 26954.2
R80 vss.n443 vss.n34 26948.4
R81 vss.n422 vss.n34 26948.4
R82 vss.n437 vss.n424 25442
R83 vss.n424 vss.n423 25442
R84 vss.n437 vss.n425 25436.2
R85 vss.n425 vss.n423 25436.2
R86 vss.n336 vss.n6 24232.3
R87 vss.n447 vss.n28 17753.2
R88 vss.n447 vss.n29 17753.2
R89 vss.n309 vss.n28 17753.2
R90 vss.n309 vss.n29 17753.2
R91 vss.n466 vss.n5 16119.1
R92 vss.n317 vss.n316 12277.7
R93 vss.n398 vss.n316 12277.7
R94 vss.n397 vss.n317 12277.7
R95 vss.n398 vss.n397 12277.7
R96 vss.n337 vss.n336 9391.71
R97 vss.n394 vss.n49 6732.77
R98 vss.n401 vss.n49 6732.77
R99 vss.n394 vss.n50 6732.77
R100 vss.n401 vss.n50 6732.77
R101 vss.n367 vss.n337 6373.53
R102 vss.n432 vss.n3 6275.03
R103 vss.n468 vss.n3 6275.03
R104 vss.n432 vss.n4 6275.03
R105 vss.n468 vss.n4 6275.03
R106 vss.n57 vss.n56 5636.95
R107 vss.n53 vss.n52 5636.95
R108 vss.n347 vss.n334 4519.41
R109 vss.n347 vss.n335 4519.41
R110 vss.n369 vss.n334 4519.41
R111 vss.n369 vss.n335 4519.41
R112 vss.n465 vss.n464 4064.84
R113 vss.n344 vss.n338 3412.74
R114 vss.n344 vss.n339 3412.74
R115 vss.n365 vss.n338 3406.94
R116 vss.n365 vss.n339 3406.94
R117 vss.n346 vss.n337 2223.62
R118 vss.n449 vss.n448 2022.67
R119 vss.n372 vss.n332 1960.4
R120 vss.n440 vss.n439 1944.26
R121 vss.t66 vss.n5 1579.6
R122 vss.n430 vss.t65 1579.6
R123 vss.n220 vss.t6 1564.71
R124 vss.n439 vss.t11 1324.96
R125 vss.n438 vss.t64 1324.96
R126 vss.n261 vss.n94 1305.6
R127 vss.n446 vss.n445 1245.36
R128 vss.n221 vss.n220 1058.82
R129 vss.n221 vss.n104 1058.82
R130 vss.n234 vss.n104 1058.82
R131 vss.n235 vss.n234 1058.82
R132 vss.n236 vss.n235 1058.82
R133 vss.n238 vss.n97 1058.82
R134 vss.n251 vss.n97 1058.82
R135 vss.n252 vss.n251 1058.82
R136 vss.n266 vss.n252 1058.82
R137 vss.n266 vss.n265 1058.82
R138 vss.n464 vss.t52 968.468
R139 vss.n265 vss.n264 951.085
R140 vss.n23 vss.n20 903.91
R141 vss.n449 vss.t52 783.348
R142 vss.n315 vss.n314 767.418
R143 vss.n236 vss.t6 717.648
R144 vss.t56 vss.n313 687.957
R145 vss.n307 vss.n306 635.574
R146 vss.n215 vss.n214 588.759
R147 vss.n218 vss.n111 588.759
R148 vss.n355 vss.n354 588.515
R149 vss.n255 vss.n96 585
R150 vss.n265 vss.n96 585
R151 vss.n268 vss.n267 585
R152 vss.n267 vss.n266 585
R153 vss.n95 vss.n93 585
R154 vss.n252 vss.n95 585
R155 vss.n250 vss.n249 585
R156 vss.n251 vss.n250 585
R157 vss.n99 vss.n98 585
R158 vss.n98 vss.n97 585
R159 vss.n240 vss.n239 585
R160 vss.n239 vss.n238 585
R161 vss.n237 vss.n102 585
R162 vss.n237 vss.n236 585
R163 vss.n107 vss.n103 585
R164 vss.n235 vss.n103 585
R165 vss.n233 vss.n232 585
R166 vss.n234 vss.n233 585
R167 vss.n224 vss.n105 585
R168 vss.n105 vss.n104 585
R169 vss.n223 vss.n222 585
R170 vss.n222 vss.n221 585
R171 vss.n219 vss.n109 585
R172 vss.n220 vss.n219 585
R173 vss.n213 vss.n117 585
R174 vss.n120 vss.n116 585
R175 vss.n217 vss.n116 585
R176 vss.n208 vss.n207 585
R177 vss.n200 vss.n123 585
R178 vss.n202 vss.n201 585
R179 vss.n193 vss.n125 585
R180 vss.n195 vss.n194 585
R181 vss.n186 vss.n182 585
R182 vss.n188 vss.n187 585
R183 vss.n184 vss.n110 585
R184 vss.n218 vss.n217 585
R185 vss.n254 vss.n253 585
R186 vss.n258 vss.n257 585
R187 vss.n83 vss.n81 585
R188 vss.n256 vss.n81 585
R189 vss.n276 vss.n275 585
R190 vss.n277 vss.n276 585
R191 vss.n87 vss.n79 585
R192 vss.n280 vss.n79 585
R193 vss.n282 vss.n80 585
R194 vss.n282 vss.n281 585
R195 vss.n287 vss.n286 585
R196 vss.n286 vss.n285 585
R197 vss.n78 vss.n76 585
R198 vss.n284 vss.n78 585
R199 vss.n72 vss.n69 585
R200 vss.n283 vss.n69 585
R201 vss.n295 vss.n294 585
R202 vss.n296 vss.n295 585
R203 vss.n70 vss.n68 585
R204 vss.n297 vss.n68 585
R205 vss.n299 vss.n60 585
R206 vss.n299 vss.n298 585
R207 vss.n263 vss.n262 585
R208 vss.n264 vss.n263 585
R209 vss.n301 vss.n300 585
R210 vss.n304 vss.n303 585
R211 vss.n143 vss.n62 585
R212 vss.n150 vss.n149 585
R213 vss.n148 vss.n142 585
R214 vss.n175 vss.n174 585
R215 vss.n173 vss.n172 585
R216 vss.n164 vss.n140 585
R217 vss.n166 vss.n165 585
R218 vss.n162 vss.n161 585
R219 vss.n160 vss.n159 585
R220 vss.n119 vss.n118 585
R221 vss.n448 vss.t46 576.794
R222 vss.n314 vss.t56 522.764
R223 vss.n355 vss.n353 512.625
R224 vss.t49 vss.t46 502.747
R225 vss.t50 vss.t49 502.747
R226 vss.t47 vss.t50 502.747
R227 vss.n431 vss.t35 493.086
R228 vss.n467 vss.t35 493.086
R229 vss.n264 vss.n253 435.913
R230 vss.n298 vss.n297 408.67
R231 vss.n297 vss.n296 408.67
R232 vss.n284 vss.n283 408.67
R233 vss.n285 vss.n284 408.67
R234 vss.n281 vss.n280 408.67
R235 vss.n257 vss.n256 408.67
R236 vss.n257 vss.n253 408.67
R237 vss.n431 vss.n430 391.663
R238 vss.n238 vss.t6 341.176
R239 vss.n442 vss.t6 314.589
R240 vss.n55 vss.t6 311.781
R241 vss.n436 vss.n426 307.036
R242 vss.n348 vss.n347 292.5
R243 vss.n347 vss.n346 292.5
R244 vss.n370 vss.n369 292.5
R245 vss.n369 vss.n368 292.5
R246 vss.n279 vss.t52 287.067
R247 vss.n308 vss.n30 281.336
R248 vss.n446 vss.n30 281.243
R249 vss.t5 vss.n441 279.022
R250 vss.n322 vss.n319 270.709
R251 vss.n256 vss.t6 267.906
R252 vss.n461 vss.n10 262.366
R253 vss.n226 vss.n108 258.334
R254 vss.n215 vss.n118 257.466
R255 vss.n436 vss.n435 256.805
R256 vss.n444 vss.n32 255.26
R257 vss.n217 vss.n216 254.34
R258 vss.n217 vss.n112 254.34
R259 vss.n217 vss.n113 254.34
R260 vss.n217 vss.n114 254.34
R261 vss.n217 vss.n115 254.34
R262 vss.n260 vss.n259 254.34
R263 vss.n306 vss.n59 254.34
R264 vss.n302 vss.n301 254.34
R265 vss.n301 vss.n67 254.34
R266 vss.n301 vss.n66 254.34
R267 vss.n301 vss.n65 254.34
R268 vss.n301 vss.n64 254.34
R269 vss.n301 vss.n63 254.34
R270 vss.n462 vss.n9 252.304
R271 vss.n296 vss.t6 249.743
R272 vss.n219 vss.n218 249.663
R273 vss.n368 vss.n318 232.525
R274 vss.n280 vss.n279 227.038
R275 vss.n451 vss.n27 223.468
R276 vss.n469 vss.n2 216.017
R277 vss.n281 vss.t6 213.417
R278 vss.n421 vss.n35 200.388
R279 vss.n442 vss.t54 199
R280 vss.n368 vss.n367 195.305
R281 vss.n285 vss.t6 195.254
R282 vss.n52 vss.n51 194.863
R283 vss.t9 vss.t41 191.542
R284 vss.n51 vss.t6 190.965
R285 vss.n400 vss.t51 189.031
R286 vss.n272 vss.n91 185
R287 vss.n274 vss.n273 185
R288 vss.n89 vss.n88 185
R289 vss.n86 vss.n85 185
R290 vss.n77 vss.n75 185
R291 vss.n289 vss.n288 185
R292 vss.n291 vss.n74 185
R293 vss.n293 vss.n292 185
R294 vss.n144 vss.n71 185
R295 vss.n145 vss.n61 185
R296 vss.n145 vss.t30 185
R297 vss.n147 vss.n146 185
R298 vss.n152 vss.n151 185
R299 vss.n153 vss.n139 185
R300 vss.n155 vss.n138 185
R301 vss.n171 vss.n170 185
R302 vss.n168 vss.n167 185
R303 vss.n163 vss.n156 185
R304 vss.n156 vss.t30 185
R305 vss.n158 vss.n157 185
R306 vss.n212 vss.n211 185
R307 vss.n210 vss.n209 185
R308 vss.n206 vss.n205 185
R309 vss.n204 vss.n203 185
R310 vss.n199 vss.n198 185
R311 vss.n197 vss.n196 185
R312 vss.n192 vss.n191 185
R313 vss.n190 vss.n189 185
R314 vss.n185 vss.n108 185
R315 vss.n270 vss.n269 185
R316 vss.n248 vss.n92 185
R317 vss.n247 vss.n246 185
R318 vss.n244 vss.n100 185
R319 vss.n242 vss.n241 185
R320 vss.n178 vss.n101 185
R321 vss.n231 vss.n230 185
R322 vss.n228 vss.n106 185
R323 vss.n226 vss.n225 185
R324 vss.n435 vss.n434 184.031
R325 vss.n279 vss.n277 181.631
R326 vss.n427 vss.n426 177.084
R327 vss.n117 vss.n116 175.546
R328 vss.n207 vss.n116 175.546
R329 vss.n201 vss.n200 175.546
R330 vss.n194 vss.n193 175.546
R331 vss.n187 vss.n186 175.546
R332 vss.n218 vss.n110 175.546
R333 vss.n161 vss.n160 175.546
R334 vss.n165 vss.n164 175.546
R335 vss.n174 vss.n173 175.546
R336 vss.n149 vss.n148 175.546
R337 vss.n303 vss.n62 175.546
R338 vss.n299 vss.n68 175.546
R339 vss.n295 vss.n68 175.546
R340 vss.n295 vss.n69 175.546
R341 vss.n78 vss.n69 175.546
R342 vss.n286 vss.n78 175.546
R343 vss.n286 vss.n282 175.546
R344 vss.n282 vss.n79 175.546
R345 vss.n276 vss.n79 175.546
R346 vss.n276 vss.n81 175.546
R347 vss.n258 vss.n81 175.546
R348 vss.n222 vss.n219 175.546
R349 vss.n222 vss.n105 175.546
R350 vss.n233 vss.n105 175.546
R351 vss.n233 vss.n103 175.546
R352 vss.n237 vss.n103 175.546
R353 vss.n239 vss.n237 175.546
R354 vss.n239 vss.n98 175.546
R355 vss.n250 vss.n98 175.546
R356 vss.n250 vss.n95 175.546
R357 vss.n267 vss.n95 175.546
R358 vss.n267 vss.n96 175.546
R359 vss.n263 vss.n96 175.546
R360 vss.n453 vss.n452 169.446
R361 vss.n145 vss.n144 163.333
R362 vss.n283 vss.t6 158.928
R363 vss.n302 vss.n59 152.643
R364 vss.n157 vss.n156 150
R365 vss.n168 vss.n156 150
R366 vss.n170 vss.n155 150
R367 vss.n153 vss.n152 150
R368 vss.n146 vss.n145 150
R369 vss.n211 vss.n210 150
R370 vss.n205 vss.n204 150
R371 vss.n198 vss.n197 150
R372 vss.n191 vss.n190 150
R373 vss.n230 vss.n228 150
R374 vss.n242 vss.n101 150
R375 vss.n246 vss.n244 150
R376 vss.n270 vss.n92 150
R377 vss.n292 vss.n291 150
R378 vss.n289 vss.n75 150
R379 vss.n89 vss.n85 150
R380 vss.n273 vss.n272 150
R381 vss.n348 vss.n342 149.538
R382 vss.n445 vss.n444 147.642
R383 vss.n300 vss.n299 146.287
R384 vss.t10 vss.n399 141.774
R385 vss.n277 vss.t6 140.764
R386 vss.n263 vss.n254 138.486
R387 vss.n420 vss.n36 137.462
R388 vss.n395 vss.n318 129.227
R389 vss.n342 vss.n332 126.4
R390 vss.n413 vss.n36 122.373
R391 vss.n404 vss.n46 113.549
R392 vss.t54 vss.t5 113.472
R393 vss.n441 vss.n440 111.778
R394 vss.n353 vss.n46 109.558
R395 vss.n373 vss.n331 104.918
R396 vss.n301 vss.t6 105.091
R397 vss.n298 vss.t6 104.439
R398 vss.n396 vss.t51 99.1166
R399 vss.n365 vss.n364 97.5005
R400 vss.n366 vss.n365 97.5005
R401 vss.n344 vss.n341 97.5005
R402 vss.n345 vss.n344 97.5005
R403 vss.n429 vss.n428 89.9525
R404 vss.n352 vss.t27 89.2211
R405 vss.n352 vss.t29 89.0687
R406 vss.t33 vss.t9 84.8974
R407 vss.t26 vss.n343 84.4265
R408 vss.n343 vss.t28 82.5503
R409 vss.n310 vss.n309 76.8967
R410 vss.n345 vss.t26 76.4529
R411 vss.n216 vss.n215 76.3222
R412 vss.n207 vss.n112 76.3222
R413 vss.n201 vss.n113 76.3222
R414 vss.n194 vss.n114 76.3222
R415 vss.n187 vss.n115 76.3222
R416 vss.n160 vss.n63 76.3222
R417 vss.n165 vss.n64 76.3222
R418 vss.n173 vss.n65 76.3222
R419 vss.n148 vss.n66 76.3222
R420 vss.n67 vss.n62 76.3222
R421 vss.n300 vss.n59 76.3222
R422 vss.n259 vss.n254 76.3222
R423 vss.n216 vss.n117 76.3222
R424 vss.n200 vss.n112 76.3222
R425 vss.n193 vss.n113 76.3222
R426 vss.n186 vss.n114 76.3222
R427 vss.n115 vss.n110 76.3222
R428 vss.n259 vss.n258 76.3222
R429 vss.n303 vss.n302 76.3222
R430 vss.n149 vss.n67 76.3222
R431 vss.n174 vss.n66 76.3222
R432 vss.n164 vss.n65 76.3222
R433 vss.n161 vss.n64 76.3222
R434 vss.n118 vss.n63 76.3222
R435 vss.n211 vss.n121 74.5978
R436 vss.n157 vss.n121 74.5978
R437 vss.n56 vss.n55 74.0483
R438 vss.n341 vss.n340 73.0981
R439 vss.n271 vss.n270 69.3109
R440 vss.n272 vss.n271 69.3109
R441 vss.n27 vss.n9 69.0601
R442 vss.n90 vss.t30 65.8183
R443 vss.n84 vss.t30 65.8183
R444 vss.n290 vss.t30 65.8183
R445 vss.t30 vss.n73 65.8183
R446 vss.n141 vss.t30 65.8183
R447 vss.n154 vss.t30 65.8183
R448 vss.n169 vss.t30 65.8183
R449 vss.n122 vss.t30 65.8183
R450 vss.n124 vss.t30 65.8183
R451 vss.n126 vss.t30 65.8183
R452 vss.n183 vss.t30 65.8183
R453 vss.n245 vss.t30 65.8183
R454 vss.n243 vss.t30 65.8183
R455 vss.n229 vss.t30 65.8183
R456 vss.n227 vss.t30 65.8183
R457 vss.n313 vss.t52 65.4995
R458 vss.n350 vss.n339 65.0005
R459 vss.n343 vss.n339 65.0005
R460 vss.n340 vss.n338 65.0005
R461 vss.n343 vss.n338 65.0005
R462 vss.n309 vss.n308 65.0005
R463 vss.n447 vss.n446 65.0005
R464 vss.n448 vss.n447 65.0005
R465 vss.t6 vss.t47 60.4079
R466 vss.t19 vss.t6 60.4079
R467 vss.t13 vss.t6 60.4079
R468 vss.n271 vss.t30 57.8461
R469 vss.n52 vss.t19 56.5107
R470 vss.n56 vss.t13 56.5107
R471 vss.n364 vss.n340 56.241
R472 vss.n121 vss.t30 55.2026
R473 vss.n18 vss.n13 54.0035
R474 vss.n16 vss.n14 54.0035
R475 vss.n407 vss.n43 53.9338
R476 vss.n409 vss.n42 53.9338
R477 vss.n169 vss.n168 53.3664
R478 vss.n155 vss.n154 53.3664
R479 vss.n152 vss.n141 53.3664
R480 vss.n210 vss.n122 53.3664
R481 vss.n204 vss.n124 53.3664
R482 vss.n197 vss.n126 53.3664
R483 vss.n190 vss.n183 53.3664
R484 vss.n227 vss.n226 53.3664
R485 vss.n230 vss.n229 53.3664
R486 vss.n243 vss.n242 53.3664
R487 vss.n246 vss.n245 53.3664
R488 vss.n292 vss.n73 53.3664
R489 vss.n290 vss.n289 53.3664
R490 vss.n85 vss.n84 53.3664
R491 vss.n273 vss.n90 53.3664
R492 vss.n90 vss.n89 53.3664
R493 vss.n84 vss.n75 53.3664
R494 vss.n291 vss.n290 53.3664
R495 vss.n144 vss.n73 53.3664
R496 vss.n146 vss.n141 53.3664
R497 vss.n154 vss.n153 53.3664
R498 vss.n170 vss.n169 53.3664
R499 vss.n205 vss.n122 53.3664
R500 vss.n198 vss.n124 53.3664
R501 vss.n191 vss.n126 53.3664
R502 vss.n183 vss.n108 53.3664
R503 vss.n245 vss.n92 53.3664
R504 vss.n244 vss.n243 53.3664
R505 vss.n229 vss.n101 53.3664
R506 vss.n228 vss.n227 53.3664
R507 vss.n4 vss.n1 53.1823
R508 vss.t35 vss.n4 53.1823
R509 vss.n3 vss.n2 53.1823
R510 vss.t35 vss.n3 53.1823
R511 vss.t6 vss.t48 53.1497
R512 vss.t6 vss.t0 53.1497
R513 vss.t6 vss.t4 53.1497
R514 vss.t6 vss.t1 53.1497
R515 vss.t6 vss.t2 53.1497
R516 vss.t6 vss.t20 53.1497
R517 vss.t6 vss.t18 53.1497
R518 vss.t6 vss.t21 53.1497
R519 vss.t6 vss.t22 53.1497
R520 vss.t6 vss.t14 53.1497
R521 vss.t6 vss.t16 53.1497
R522 vss.t6 vss.t12 53.1497
R523 vss.t6 vss.t15 53.1497
R524 vss.n399 vss.n315 49.7676
R525 vss.n402 vss.n401 48.7505
R526 vss.n401 vss.n400 48.7505
R527 vss.n394 vss.n393 48.7505
R528 vss.n395 vss.n394 48.7505
R529 vss.n366 vss.t24 45.4967
R530 vss.n311 vss.n310 44.185
R531 vss.n470 vss.n469 42.0571
R532 vss.n435 vss.n2 41.1681
R533 vss.n367 vss.n366 39.8683
R534 vss.n22 vss.n21 39.7638
R535 vss.n453 vss.n24 39.511
R536 vss.n278 vss.t3 39.3863
R537 vss.n342 vss.n335 34.4123
R538 vss.t24 vss.n335 34.4123
R539 vss.n351 vss.n334 34.4123
R540 vss.t24 vss.n334 34.4123
R541 vss.n469 vss.n468 34.4123
R542 vss.n468 vss.n467 34.4123
R543 vss.n433 vss.n432 34.4123
R544 vss.n432 vss.n431 34.4123
R545 vss.n404 vss.n403 33.9329
R546 vss.n326 vss.n50 32.5005
R547 vss.t33 vss.n50 32.5005
R548 vss.n375 vss.n49 32.5005
R549 vss.t33 vss.n49 32.5005
R550 vss.n22 vss.n8 32.5005
R551 vss.n440 vss.n8 32.5005
R552 vss.n27 vss.n7 32.5005
R553 vss.n314 vss.n7 32.5005
R554 vss.t28 vss.t24 32.3638
R555 vss.n421 vss.n420 32.1396
R556 vss.n1 vss.t36 30.8834
R557 vss.n363 vss.n333 30.4707
R558 vss.n346 vss.n345 28.6115
R559 vss.n326 vss.n320 28.0594
R560 vss.n130 vss.t31 26.6016
R561 vss.n37 vss.t67 25.1357
R562 vss.n376 vss.n374 24.7516
R563 vss.n403 vss.n47 24.4644
R564 vss.n445 vss.n31 23.8095
R565 vss.n308 vss.n307 23.4151
R566 vss.n428 vss.n427 23.0405
R567 vss.n135 vss.n127 20.7857
R568 vss.n134 vss.n128 20.7857
R569 vss.n130 vss.n129 20.7857
R570 vss.n411 vss.n41 20.7665
R571 vss.n412 vss.n40 20.7665
R572 vss.n415 vss.n39 20.7665
R573 vss.n416 vss.n38 20.7665
R574 vss.n349 vss.n348 20.517
R575 vss.n397 vss.n47 20.1729
R576 vss.n397 vss.n396 20.1729
R577 vss.n356 vss.n316 20.1729
R578 vss.n396 vss.n316 20.1729
R579 vss.n349 vss.n341 20.0772
R580 vss.n388 vss.n387 19.4026
R581 vss.t41 vss.n395 19.2382
R582 vss.n392 vss.n320 19.2005
R583 vss.n398 vss.n46 18.8715
R584 vss.n399 vss.n398 18.8715
R585 vss.n354 vss.n317 18.8715
R586 vss.n318 vss.n317 18.8715
R587 vss.n433 vss.n429 18.7337
R588 vss.n307 vss.n58 17.5097
R589 vss.n374 vss.n319 17.1218
R590 vss.n387 vss.n48 16.4046
R591 vss.n434 vss.n433 16.3845
R592 vss.n403 vss.n402 16.1396
R593 vss.n132 vss.n131 16.0068
R594 vss.n462 vss.n461 15.5385
R595 vss.n422 vss.n421 14.6255
R596 vss.n442 vss.n422 14.6255
R597 vss.n444 vss.n443 14.6255
R598 vss.n443 vss.n442 14.6255
R599 vss.n329 vss.n328 14.0913
R600 vss.n387 vss.n386 12.7191
R601 vss.n279 vss.n278 12.1537
R602 vss.n434 vss.n425 11.9393
R603 vss.n430 vss.n425 11.9393
R604 vss.n426 vss.n424 11.9393
R605 vss.n424 vss.n5 11.9393
R606 vss.n43 vss.t61 11.6005
R607 vss.n43 vss.t58 11.6005
R608 vss.n42 vss.t53 11.6005
R609 vss.n42 vss.t55 11.6005
R610 vss.n13 vss.t59 11.6005
R611 vss.n13 vss.t60 11.6005
R612 vss.n14 vss.t57 11.6005
R613 vss.n14 vss.t62 11.6005
R614 vss.n452 vss.n451 10.5495
R615 vss.n429 vss.n1 10.0532
R616 vss.n371 vss.n333 9.74099
R617 vss.n390 vss.n322 9.3005
R618 vss.n454 vss.n453 9.3005
R619 vss.n459 vss.n10 9.3005
R620 vss.n20 vss.n12 9.3005
R621 vss.n350 vss.n349 8.86924
R622 vss.n370 vss.n332 8.42977
R623 vss.n396 vss.t33 7.5283
R624 vss.n427 vss.n423 7.5005
R625 vss.n438 vss.n423 7.5005
R626 vss.n437 vss.n436 7.5005
R627 vss.n438 vss.n437 7.5005
R628 vss.n376 vss.n375 7.34725
R629 vss.n373 vss.n372 7.32557
R630 vss.n31 vss.n29 7.313
R631 vss.n51 vss.n29 7.313
R632 vss.n30 vss.n28 7.313
R633 vss.n51 vss.n28 7.313
R634 vss.n374 vss.n373 6.9983
R635 vss.n420 vss.n419 6.9005
R636 vss.n418 vss.n36 6.9005
R637 vss.n385 vss 6.21282
R638 vss.n58 vss.n33 6.15839
R639 vss.n55 vss.n33 6.15839
R640 vss.n34 vss.n32 6.15839
R641 vss.n441 vss.n34 6.15839
R642 vss.n363 vss.n362 5.92892
R643 vss.n372 vss.n371 5.77749
R644 vss.n351 vss.n350 5.73359
R645 vss.n364 vss.n363 5.34506
R646 vss.n278 vss.t6 4.95804
R647 vss.n159 vss.n119 4.90263
R648 vss.n223 vss.n109 4.90263
R649 vss.n451 vss.n450 4.8755
R650 vss.n450 vss.n449 4.8755
R651 vss.n463 vss.n462 4.8755
R652 vss.n464 vss.n463 4.8755
R653 vss.n225 vss.n223 4.84816
R654 vss.n224 vss.n106 4.84816
R655 vss.n232 vss.n231 4.84816
R656 vss.n241 vss.n102 4.84816
R657 vss.n240 vss.n100 4.84816
R658 vss.n247 vss.n99 4.84816
R659 vss.n249 vss.n248 4.84816
R660 vss.n269 vss.n93 4.84816
R661 vss.n262 vss.n255 4.57193
R662 vss.n454 vss.n26 4.5005
R663 vss.n386 vss.n385 4.5005
R664 vss.n45 vss.n44 4.5005
R665 vss.n390 vss.n323 4.5005
R666 vss.n459 vss.n458 4.5005
R667 vss.n457 vss.n12 4.5005
R668 vss.n41 vss.t32 4.3505
R669 vss.n41 vss.t7 4.3505
R670 vss.n40 vss.t44 4.3505
R671 vss.n40 vss.t23 4.3505
R672 vss.n39 vss.t45 4.3505
R673 vss.n39 vss.t38 4.3505
R674 vss.n38 vss.t42 4.3505
R675 vss.n38 vss.t25 4.3505
R676 vss.n127 vss.t63 4.3505
R677 vss.n127 vss.t40 4.3505
R678 vss.n128 vss.t8 4.3505
R679 vss.n128 vss.t17 4.3505
R680 vss.n129 vss.t43 4.3505
R681 vss.n129 vss.t39 4.3505
R682 vss.n457 vss.n0 4.26937
R683 vss.n15 vss.n11 4.25229
R684 vss.n460 vss.n459 4.1668
R685 vss.n419 vss.n37 4.10351
R686 vss.n16 vss.n15 4.02718
R687 vss.n407 vss.n406 3.98965
R688 vss.n354 vss.n331 3.98739
R689 vss.n260 vss.n35 3.9624
R690 vss.n159 vss.n158 3.81327
R691 vss.n163 vss.n162 3.81327
R692 vss.n167 vss.n166 3.81327
R693 vss.n171 vss.n140 3.81327
R694 vss.n172 vss.n138 3.81327
R695 vss.n175 vss.n139 3.81327
R696 vss.n151 vss.n142 3.81327
R697 vss.n150 vss.n147 3.81327
R698 vss.n143 vss.n61 3.81327
R699 vss.n21 vss.n10 3.76521
R700 vss.n470 vss.n1 3.71562
R701 vss.n255 vss.n94 3.55606
R702 vss.n179 vss.n178 3.48646
R703 vss.n471 vss.n0 3.33015
R704 vss.n328 vss.t37 3.16414
R705 vss.n328 vss.t34 3.16414
R706 vss.n15 vss.n9 3.10035
R707 vss.n388 vss.n326 2.96471
R708 vss.n217 vss.t6 128.062
R709 vss.n213 vss.n212 2.7239
R710 vss.n209 vss.n120 2.7239
R711 vss.n208 vss.n206 2.7239
R712 vss.n203 vss.n123 2.7239
R713 vss.n202 vss.n199 2.7239
R714 vss.n195 vss.n192 2.7239
R715 vss.n189 vss.n182 2.7239
R716 vss.n188 vss.n185 2.7239
R717 vss.n358 vss.n357 2.68591
R718 vss.n400 vss.t10 2.50977
R719 vss.n360 vss.n333 2.3255
R720 vss.n454 vss.n25 2.29617
R721 vss.n419 vss.n418 2.28754
R722 vss.n456 vss.n19 2.24795
R723 vss.n212 vss.n120 2.17922
R724 vss.n209 vss.n208 2.17922
R725 vss.n206 vss.n123 2.17922
R726 vss.n203 vss.n202 2.17922
R727 vss.n199 vss.n125 2.17922
R728 vss.n196 vss.n195 2.17922
R729 vss.n192 vss.n182 2.17922
R730 vss.n189 vss.n188 2.17922
R731 vss.n185 vss.n184 2.17922
R732 vss.n70 vss.n60 2.17819
R733 vss.n17 vss.n16 2.15904
R734 vss.n458 vss.n18 2.12067
R735 vss.n357 vss.n353 2.10102
R736 vss.n136 vss.n82 1.89157
R737 vss.n294 vss.n71 1.79105
R738 vss.n293 vss.n72 1.79105
R739 vss.n76 vss.n74 1.79105
R740 vss.n288 vss.n287 1.79105
R741 vss.n80 vss.n77 1.79105
R742 vss.n274 vss.n83 1.79105
R743 vss.n18 vss.n17 1.78099
R744 vss.n471 vss.n470 1.7255
R745 vss.n131 vss 1.7155
R746 vss.n181 vss.n125 1.68901
R747 vss.n411 vss.n410 1.67152
R748 vss.n306 vss.n305 1.64587
R749 vss.n312 vss.t6 1.63432
R750 vss.n359 vss.n358 1.55732
R751 vss.n180 vss.n179 1.51978
R752 vss.n362 vss.n351 1.47378
R753 vss.n135 vss.n134 1.46641
R754 vss.n133 vss.n130 1.43989
R755 vss.n87 vss 1.37971
R756 vss.n91 vss.n35 1.37971
R757 vss.n310 vss.t6 1.37561
R758 vss.n179 vss.n107 1.3622
R759 vss.n24 vss.n23 1.30961
R760 vss.n408 vss.n407 1.23783
R761 vss.n275 vss.n82 1.18613
R762 vss.n410 vss.n409 1.13184
R763 vss.n261 vss.n260 1.11796
R764 vss.n162 vss.n158 1.08986
R765 vss.n166 vss.n163 1.08986
R766 vss.n167 vss.n140 1.08986
R767 vss.n172 vss.n171 1.08986
R768 vss.n142 vss.n139 1.08986
R769 vss.n151 vss.n150 1.08986
R770 vss.n147 vss.n143 1.08986
R771 vss.n304 vss.n61 1.08986
R772 vss.n305 vss.n304 1.08986
R773 vss.n268 vss.n94 1.08986
R774 vss.t11 vss.t66 1.07946
R775 vss.n439 vss.n438 1.07946
R776 vss.t65 vss.t64 1.07946
R777 vss.n406 vss.n44 1.07186
R778 vss.n23 vss.n22 1.06085
R779 vss.n405 vss.n45 1.05279
R780 vss.n196 vss.n181 1.03539
R781 vss.n405 vss.n404 1.03383
R782 vss.n412 vss.n411 0.998567
R783 vss.n416 vss.n415 0.997923
R784 vss.n409 vss.n408 0.995892
R785 vss.n176 vss.n138 0.871989
R786 vss.n214 vss.n119 0.817521
R787 vss.n111 vss.n109 0.817521
R788 vss.n305 vss.n60 0.798988
R789 vss.n322 vss.n320 0.775237
R790 vss.n180 vss.n177 0.765632
R791 vss.n132 vss.n58 0.739443
R792 vss.n21 vss.n20 0.684992
R793 vss.n375 vss.n47 0.682157
R794 vss.n177 vss.n137 0.653909
R795 vss.n417 vss.n416 0.633876
R796 vss.n88 vss.n82 0.605415
R797 vss.n181 vss.n180 0.596304
R798 vss.n177 vss.n176 0.59175
R799 vss.n137 vss.n135 0.539326
R800 vss.n413 vss.n32 0.532356
R801 vss.n414 vss.n412 0.528206
R802 vss.n390 vss.n389 0.47062
R803 vss.n415 vss.n414 0.469572
R804 vss.n455 vss.n454 0.469344
R805 vss.n324 vss.n323 0.456098
R806 vss.n137 vss.n136 0.452967
R807 vss.n379 vss.n377 0.452003
R808 vss.n406 vss.n405 0.4505
R809 vss.n455 vss.n12 0.441368
R810 vss vss.n86 0.411842
R811 vss.n323 vss.n321 0.399345
R812 vss.n357 vss.n356 0.391918
R813 vss.n71 vss.n70 0.387646
R814 vss.n294 vss.n293 0.387646
R815 vss.n74 vss.n72 0.387646
R816 vss.n288 vss.n76 0.387646
R817 vss.n287 vss.n77 0.387646
R818 vss.n88 vss.n87 0.387646
R819 vss.n275 vss.n274 0.387646
R820 vss.n91 vss.n83 0.387646
R821 vss.n377 vss.n330 0.376108
R822 vss.n360 vss.n359 0.368932
R823 vss.n361 vss.n360 0.355
R824 vss.n389 vss.n325 0.350102
R825 vss.n327 vss.n324 0.344129
R826 vss.n418 vss.n417 0.343093
R827 vss.n455 vss.n24 0.32741
R828 vss.n214 vss.n213 0.327309
R829 vss.n379 vss.n378 0.326722
R830 vss.n457 vss.n456 0.317677
R831 vss.n330 vss.n321 0.312188
R832 vss.n358 vss.n331 0.3005
R833 vss.n391 vss.n390 0.272145
R834 vss vss.n80 0.242466
R835 vss.n384 vss.n383 0.226831
R836 vss.n393 vss.n319 0.224276
R837 vss.n392 vss.n391 0.221929
R838 vss.n380 vss.n379 0.221128
R839 vss.n382 vss.n325 0.220839
R840 vss.n176 vss.n175 0.218372
R841 vss.n378 vss.n329 0.216846
R842 vss.n381 vss.n380 0.20954
R843 vss.n131 vss.n31 0.188367
R844 vss.n371 vss.n370 0.187817
R845 vss.n356 vss.n355 0.180782
R846 vss.n86 vss 0.14568
R847 vss.n428 vss.n0 0.139042
R848 vss.n381 vss.n48 0.133357
R849 vss.n377 vss.n376 0.126176
R850 vss.n456 vss.n455 0.1255
R851 vss.n362 vss.n361 0.122868
R852 vss vss.n471 0.120187
R853 vss.n361 vss.n352 0.118284
R854 vss.n184 vss.n111 0.109436
R855 vss.n389 vss.n388 0.107397
R856 vss.n133 vss.n132 0.0987955
R857 vss.n136 vss.n37 0.0948141
R858 vss.n19 vss 0.0874816
R859 vss.n410 vss.n26 0.0851774
R860 vss.n461 vss.n460 0.0850455
R861 vss.n417 vss 0.0849072
R862 vss.n414 vss.n413 0.0736577
R863 vss.n459 vss.n12 0.0711522
R864 vss.n383 vss.n382 0.0605
R865 vss.n225 vss.n224 0.0549681
R866 vss.n232 vss.n106 0.0549681
R867 vss.n231 vss.n107 0.0549681
R868 vss.n178 vss.n102 0.0549681
R869 vss.n241 vss.n240 0.0549681
R870 vss.n100 vss.n99 0.0549681
R871 vss.n249 vss.n247 0.0549681
R872 vss.n248 vss.n93 0.0549681
R873 vss.n269 vss.n268 0.0549681
R874 vss.n262 vss.n261 0.0512937
R875 vss vss.n384 0.048119
R876 vss.n389 vss.n324 0.0459545
R877 vss.n393 vss.n392 0.0452552
R878 vss.n385 vss.n327 0.0448787
R879 vss.n386 vss.n325 0.0428729
R880 vss.n359 vss.n330 0.0382747
R881 vss.n17 vss.n11 0.0367903
R882 vss.n378 vss.n44 0.0330444
R883 vss.n380 vss.n45 0.0294548
R884 vss.n452 vss.n25 0.0286818
R885 vss.n134 vss.n133 0.0270152
R886 vss.n402 vss.n48 0.027001
R887 vss.n458 vss.n457 0.0246098
R888 vss.n26 vss.n19 0.0195092
R889 vss.n460 vss.n11 0.0135435
R890 vss.n408 vss.n25 0.0126951
R891 vss.n391 vss.n321 0.00969913
R892 vss.n384 vss.n327 0.00493787
R893 vss.n383 vss.n329 0.00234911
R894 vss.n382 vss.n381 0.00191243
R895 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 935.75
R896 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 235.982
R897 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 235.978
R898 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 190.305
R899 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 190.305
R900 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 190.305
R901 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 190.305
R902 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 190.305
R903 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 190.305
R904 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 95.3928
R905 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 95.3648
R906 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 95.1789
R907 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 95.1648
R908 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 95.1542
R909 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 95.1535
R910 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 94.8314
R911 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 94.8314
R912 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 94.8314
R913 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 94.8314
R914 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 94.8314
R915 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 94.8314
R916 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 94.8314
R917 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 94.8314
R918 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 94.8314
R919 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 94.8314
R920 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 94.8314
R921 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 94.8314
R922 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 94.8314
R923 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 94.8314
R924 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 94.8314
R925 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 94.8314
R926 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 94.8314
R927 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 94.8314
R928 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 94.8314
R929 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 94.8314
R930 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 94.8314
R931 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 94.8314
R932 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 94.8314
R933 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 84.0884
R934 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 83.5719
R935 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 83.5719
R936 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 83.5719
R937 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 83.5719
R938 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 73.19
R939 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 26.074
R940 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 26.074
R941 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 26.074
R942 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 25.7843
R943 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 10.2822
R944 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 9.66398
R945 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R946 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R947 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R948 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R949 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R950 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 9.3005
R951 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R952 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R953 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 9.3005
R954 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R955 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R956 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R957 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R958 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R959 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R960 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R961 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R962 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R963 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R964 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R965 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R966 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R967 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 9.3005
R968 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R969 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R970 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 9.3005
R971 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 9.3005
R972 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 9.3005
R973 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 7.22993
R974 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 7.22993
R975 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 7.22993
R976 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 6.83022
R977 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 6.81633
R978 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 6.81633
R979 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 6.81633
R980 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 6.75312
R981 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 4.64588
R982 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 4.64588
R983 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 4.64588
R984 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 4.64588
R985 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 2.29815
R986 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 1.86108
R987 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 1.86108
R988 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 1.86108
R989 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 1.86108
R990 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 1.86108
R991 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 1.86108
R992 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 1.86108
R993 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 1.28692
R994 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 1.25468
R995 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 1.14402
R996 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 1.1424
R997 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 1.12066
R998 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 1.12066
R999 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 1.11251
R1000 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 1.10979
R1001 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 1.10164
R1002 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 1.10164
R1003 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 1.10164
R1004 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 1.10164
R1005 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 1.09892
R1006 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 1.09349
R1007 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 1.09349
R1008 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 1.08805
R1009 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 1.08262
R1010 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 1.08262
R1011 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 1.08262
R1012 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 1.07024
R1013 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 1.0237
R1014 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.959578
R1015 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 0.812055
R1016 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.77514
R1017 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.701365
R1018 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.645119
R1019 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 0.645119
R1020 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 0.645119
R1021 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 0.645119
R1022 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 0.645119
R1023 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 0.645119
R1024 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 0.645119
R1025 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.645119
R1026 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 0.645119
R1027 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.645119
R1028 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 0.645119
R1029 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 0.645119
R1030 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 0.645119
R1031 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 0.645119
R1032 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 0.645119
R1033 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.645119
R1034 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 0.645119
R1035 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.645119
R1036 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 0.645119
R1037 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 0.645119
R1038 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 0.645119
R1039 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 0.645119
R1040 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 0.645119
R1041 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.645119
R1042 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.645119
R1043 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 0.645119
R1044 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 0.645119
R1045 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 0.645119
R1046 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 0.645119
R1047 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 0.645118
R1048 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 0.590702
R1049 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 0.572258
R1050 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 0.495065
R1051 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.495065
R1052 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 0.481478
R1053 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.481478
R1054 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.475521
R1055 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 0.470609
R1056 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.470609
R1057 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 0.465174
R1058 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 0.465174
R1059 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.465174
R1060 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.459844
R1061 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 0.459739
R1062 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.459739
R1063 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 0.446152
R1064 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.446152
R1065 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.445943
R1066 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.443435
R1067 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.440717
R1068 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 0.440717
R1069 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.434551
R1070 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 0.432263
R1071 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.414484
R1072 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.408265
R1073 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.408265
R1074 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.40372
R1075 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.40372
R1076 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.314045
R1077 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 0.290206
R1078 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.0183279
R1079 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 0.0112346
R1080 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 0.0112346
R1081 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 0.0112346
R1082 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 0.0112346
R1083 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.0112346
R1084 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 0.0112346
R1085 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 0.0112346
R1086 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 0.0112346
R1087 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 0.00759293
R1088 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 0.00316393
R1089 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.t0 88.7532
R1090 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 22.2005
R1091 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 21.8665
R1092 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 21.5445
R1093 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 21.5445
R1094 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 21.5445
R1095 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 21.5445
R1096 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 21.5445
R1097 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 21.5445
R1098 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 21.5445
R1099 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 21.5445
R1100 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 21.5445
R1101 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 21.5445
R1102 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 21.5445
R1103 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 21.5445
R1104 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 21.5445
R1105 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 21.5418
R1106 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 4.3505
R1107 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 4.3505
R1108 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 4.3505
R1109 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 4.3505
R1110 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 4.3505
R1111 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 4.3505
R1112 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 4.3505
R1113 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 4.3505
R1114 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 4.3505
R1115 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 4.3505
R1116 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 4.3505
R1117 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 4.3505
R1118 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 4.3505
R1119 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 4.3505
R1120 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 4.3505
R1121 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 4.3505
R1122 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 4.3505
R1123 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 4.3505
R1124 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 4.3505
R1125 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 4.3505
R1126 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 4.3505
R1127 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 4.3505
R1128 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 4.3505
R1129 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 4.3505
R1130 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 OTA_vref_0.OTA_vref_stage2_0.vref0.t32 4.3505
R1131 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 4.3505
R1132 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 4.3505
R1133 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 4.3505
R1134 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 4.3505
R1135 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 4.3505
R1136 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 4.3505
R1137 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 4.3505
R1138 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 4.27517
R1139 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 3.08331
R1140 a_n1236_n9479.n58 a_n1236_n9479.t8 190.305
R1141 a_n1236_n9479.t8 a_n1236_n9479.n57 190.305
R1142 a_n1236_n9479.t26 a_n1236_n9479.n42 190.305
R1143 a_n1236_n9479.n56 a_n1236_n9479.t26 190.305
R1144 a_n1236_n9479.n23 a_n1236_n9479.t16 190.305
R1145 a_n1236_n9479.n21 a_n1236_n9479.t16 190.305
R1146 a_n1236_n9479.t30 a_n1236_n9479.n18 190.305
R1147 a_n1236_n9479.n20 a_n1236_n9479.t30 190.305
R1148 a_n1236_n9479.t12 a_n1236_n9479.n77 190.305
R1149 a_n1236_n9479.n81 a_n1236_n9479.t12 190.305
R1150 a_n1236_n9479.t22 a_n1236_n9479.n79 190.305
R1151 a_n1236_n9479.n80 a_n1236_n9479.t22 190.305
R1152 a_n1236_n9479.t10 a_n1236_n9479.n47 190.305
R1153 a_n1236_n9479.n48 a_n1236_n9479.t10 190.305
R1154 a_n1236_n9479.t24 a_n1236_n9479.n45 190.305
R1155 a_n1236_n9479.n49 a_n1236_n9479.t24 190.305
R1156 a_n1236_n9479.t28 a_n1236_n9479.n28 190.305
R1157 a_n1236_n9479.n32 a_n1236_n9479.t28 190.305
R1158 a_n1236_n9479.t2 a_n1236_n9479.n30 190.305
R1159 a_n1236_n9479.n31 a_n1236_n9479.t2 190.305
R1160 a_n1236_n9479.t18 a_n1236_n9479.n70 190.305
R1161 a_n1236_n9479.n71 a_n1236_n9479.t18 190.305
R1162 a_n1236_n9479.n16 a_n1236_n9479.t6 190.305
R1163 a_n1236_n9479.t6 a_n1236_n9479.n13 190.305
R1164 a_n1236_n9479.t20 a_n1236_n9479.n62 190.305
R1165 a_n1236_n9479.n63 a_n1236_n9479.t20 190.305
R1166 a_n1236_n9479.t4 a_n1236_n9479.n37 190.305
R1167 a_n1236_n9479.n64 a_n1236_n9479.t4 190.305
R1168 a_n1236_n9479.n25 a_n1236_n9479.t14 95.1811
R1169 a_n1236_n9479.n41 a_n1236_n9479.t0 95.1783
R1170 a_n1236_n9479.n54 a_n1236_n9479.n53 22.3176
R1171 a_n1236_n9479.n36 a_n1236_n9479.n35 22.2301
R1172 a_n1236_n9479.n9 a_n1236_n9479.n26 22.2284
R1173 a_n1236_n9479.n0 a_n1236_n9479.n27 22.2284
R1174 a_n1236_n9479.n6 a_n1236_n9479.n34 22.2284
R1175 a_n1236_n9479.n12 a_n1236_n9479.n69 22.2284
R1176 a_n1236_n9479.n68 a_n1236_n9479.n67 22.2284
R1177 a_n1236_n9479.n10 a_n1236_n9479.n38 22.2284
R1178 a_n1236_n9479.n40 a_n1236_n9479.n39 22.2284
R1179 a_n1236_n9479.n5 a_n1236_n9479.n17 22.1884
R1180 a_n1236_n9479.n1 a_n1236_n9479.n83 22.1884
R1181 a_n1236_n9479.n3 a_n1236_n9479.n43 22.1884
R1182 a_n1236_n9479.n2 a_n1236_n9479.n44 22.1884
R1183 a_n1236_n9479.n11 a_n1236_n9479.n51 22.1884
R1184 a_n1236_n9479.n8 a_n1236_n9479.n52 22.1884
R1185 a_n1236_n9479.n84 a_n1236_n9479.n4 22.1884
R1186 a_n1236_n9479.n59 a_n1236_n9479.n41 11.5566
R1187 a_n1236_n9479.n25 a_n1236_n9479.n24 10.9335
R1188 a_n1236_n9479.n77 a_n1236_n9479.n76 9.89233
R1189 a_n1236_n9479.n47 a_n1236_n9479.n15 9.89233
R1190 a_n1236_n9479.n24 a_n1236_n9479.n23 9.80925
R1191 a_n1236_n9479.n59 a_n1236_n9479.n58 9.80925
R1192 a_n1236_n9479.n64 a_n1236_n9479.n60 9.48127
R1193 a_n1236_n9479.n75 a_n1236_n9479.n13 9.40378
R1194 a_n1236_n9479.n31 a_n1236_n9479.n14 9.39819
R1195 a_n1236_n9479.n41 a_n1236_n9479.n40 4.9275
R1196 a_n1236_n9479.n9 a_n1236_n9479.n25 4.79654
R1197 a_n1236_n9479.n61 a_n1236_n9479.n10 4.5005
R1198 a_n1236_n9479.n66 a_n1236_n9479.n65 4.5005
R1199 a_n1236_n9479.n12 a_n1236_n9479.n72 4.5005
R1200 a_n1236_n9479.n74 a_n1236_n9479.n73 4.5005
R1201 a_n1236_n9479.n6 a_n1236_n9479.n33 4.5005
R1202 a_n1236_n9479.n29 a_n1236_n9479.n0 4.5005
R1203 a_n1236_n9479.n8 a_n1236_n9479.n7 4.5005
R1204 a_n1236_n9479.n55 a_n1236_n9479.n54 4.5005
R1205 a_n1236_n9479.n11 a_n1236_n9479.n50 4.5005
R1206 a_n1236_n9479.n46 a_n1236_n9479.n2 4.5005
R1207 a_n1236_n9479.n78 a_n1236_n9479.n3 4.5005
R1208 a_n1236_n9479.n1 a_n1236_n9479.n82 4.5005
R1209 a_n1236_n9479.n22 a_n1236_n9479.n5 4.5005
R1210 a_n1236_n9479.n19 a_n1236_n9479.n4 4.5005
R1211 a_n1236_n9479.n17 a_n1236_n9479.t37 4.3505
R1212 a_n1236_n9479.n17 a_n1236_n9479.t17 4.3505
R1213 a_n1236_n9479.n83 a_n1236_n9479.t35 4.3505
R1214 a_n1236_n9479.n83 a_n1236_n9479.t13 4.3505
R1215 a_n1236_n9479.n43 a_n1236_n9479.t23 4.3505
R1216 a_n1236_n9479.n43 a_n1236_n9479.t47 4.3505
R1217 a_n1236_n9479.n44 a_n1236_n9479.t34 4.3505
R1218 a_n1236_n9479.n44 a_n1236_n9479.t11 4.3505
R1219 a_n1236_n9479.n51 a_n1236_n9479.t25 4.3505
R1220 a_n1236_n9479.n51 a_n1236_n9479.t32 4.3505
R1221 a_n1236_n9479.n52 a_n1236_n9479.t43 4.3505
R1222 a_n1236_n9479.n52 a_n1236_n9479.t9 4.3505
R1223 a_n1236_n9479.n26 a_n1236_n9479.t15 4.3505
R1224 a_n1236_n9479.n26 a_n1236_n9479.t36 4.3505
R1225 a_n1236_n9479.n27 a_n1236_n9479.t39 4.3505
R1226 a_n1236_n9479.n27 a_n1236_n9479.t3 4.3505
R1227 a_n1236_n9479.n34 a_n1236_n9479.t29 4.3505
R1228 a_n1236_n9479.n34 a_n1236_n9479.t45 4.3505
R1229 a_n1236_n9479.n35 a_n1236_n9479.t40 4.3505
R1230 a_n1236_n9479.n35 a_n1236_n9479.t7 4.3505
R1231 a_n1236_n9479.n69 a_n1236_n9479.t19 4.3505
R1232 a_n1236_n9479.n69 a_n1236_n9479.t44 4.3505
R1233 a_n1236_n9479.n67 a_n1236_n9479.t41 4.3505
R1234 a_n1236_n9479.n67 a_n1236_n9479.t5 4.3505
R1235 a_n1236_n9479.n38 a_n1236_n9479.t21 4.3505
R1236 a_n1236_n9479.n38 a_n1236_n9479.t38 4.3505
R1237 a_n1236_n9479.n39 a_n1236_n9479.t42 4.3505
R1238 a_n1236_n9479.n39 a_n1236_n9479.t1 4.3505
R1239 a_n1236_n9479.n53 a_n1236_n9479.t27 4.3505
R1240 a_n1236_n9479.n53 a_n1236_n9479.t33 4.3505
R1241 a_n1236_n9479.t31 a_n1236_n9479.n84 4.3505
R1242 a_n1236_n9479.n84 a_n1236_n9479.t46 4.3505
R1243 a_n1236_n9479.n9 a_n1236_n9479.n5 2.55258
R1244 a_n1236_n9479.n24 a_n1236_n9479.n14 1.86108
R1245 a_n1236_n9479.n76 a_n1236_n9479.n14 1.86108
R1246 a_n1236_n9479.n76 a_n1236_n9479.n75 1.86108
R1247 a_n1236_n9479.n75 a_n1236_n9479.n15 1.86108
R1248 a_n1236_n9479.n60 a_n1236_n9479.n15 1.86108
R1249 a_n1236_n9479.n60 a_n1236_n9479.n59 1.86108
R1250 a_n1236_n9479.n0 a_n1236_n9479.n9 1.20675
R1251 a_n1236_n9479.n36 a_n1236_n9479.n6 1.0755
R1252 a_n1236_n9479.n12 a_n1236_n9479.n68 1.0755
R1253 a_n1236_n9479.n40 a_n1236_n9479.n10 1.0755
R1254 a_n1236_n9479.n8 a_n1236_n9479.n11 1.0755
R1255 a_n1236_n9479.n2 a_n1236_n9479.n3 1.0755
R1256 a_n1236_n9479.n4 a_n1236_n9479.n1 1.0755
R1257 a_n1236_n9479.n72 a_n1236_n9479.n70 0.759759
R1258 a_n1236_n9479.n74 a_n1236_n9479.n16 0.756673
R1259 a_n1236_n9479.n65 a_n1236_n9479.n37 0.702205
R1260 a_n1236_n9479.n62 a_n1236_n9479.n61 0.700784
R1261 a_n1236_n9479.n80 a_n1236_n9479.n78 0.669534
R1262 a_n1236_n9479.n48 a_n1236_n9479.n46 0.668114
R1263 a_n1236_n9479.n57 a_n1236_n9479.n7 0.666693
R1264 a_n1236_n9479.n82 a_n1236_n9479.n81 0.665273
R1265 a_n1236_n9479.n20 a_n1236_n9479.n19 0.662432
R1266 a_n1236_n9479.n22 a_n1236_n9479.n21 0.661011
R1267 a_n1236_n9479.n56 a_n1236_n9479.n55 0.659208
R1268 a_n1236_n9479.n13 a_n1236_n9479.n74 0.647608
R1269 a_n1236_n9479.n72 a_n1236_n9479.n71 0.645562
R1270 a_n1236_n9479.n23 a_n1236_n9479.n22 0.632599
R1271 a_n1236_n9479.n19 a_n1236_n9479.n18 0.631182
R1272 a_n1236_n9479.n50 a_n1236_n9479.n49 0.629532
R1273 a_n1236_n9479.n82 a_n1236_n9479.n77 0.628338
R1274 a_n1236_n9479.n58 a_n1236_n9479.n7 0.626917
R1275 a_n1236_n9479.n47 a_n1236_n9479.n46 0.625497
R1276 a_n1236_n9479.n79 a_n1236_n9479.n78 0.62408
R1277 a_n1236_n9479.n55 a_n1236_n9479.n42 0.619882
R1278 a_n1236_n9479.n50 a_n1236_n9479.n45 0.594586
R1279 a_n1236_n9479.n63 a_n1236_n9479.n61 0.59283
R1280 a_n1236_n9479.n65 a_n1236_n9479.n64 0.591408
R1281 a_n1236_n9479.n30 a_n1236_n9479.n29 0.580689
R1282 a_n1236_n9479.n33 a_n1236_n9479.n28 0.57833
R1283 a_n1236_n9479.n5 a_n1236_n9479.n4 0.538
R1284 a_n1236_n9479.n6 a_n1236_n9479.n0 0.538
R1285 a_n1236_n9479.n11 a_n1236_n9479.n2 0.537105
R1286 a_n1236_n9479.n1 a_n1236_n9479.n3 0.536664
R1287 a_n1236_n9479.n33 a_n1236_n9479.n32 0.495783
R1288 a_n1236_n9479.n31 a_n1236_n9479.n29 0.493424
R1289 a_n1236_n9479.n71 a_n1236_n9479.n13 0.488952
R1290 a_n1236_n9479.n70 a_n1236_n9479.n16 0.486913
R1291 a_n1236_n9479.n58 a_n1236_n9479.n42 0.476043
R1292 a_n1236_n9479.n57 a_n1236_n9479.n56 0.476043
R1293 a_n1236_n9479.n23 a_n1236_n9479.n18 0.459739
R1294 a_n1236_n9479.n21 a_n1236_n9479.n20 0.459739
R1295 a_n1236_n9479.n79 a_n1236_n9479.n77 0.459739
R1296 a_n1236_n9479.n81 a_n1236_n9479.n80 0.459739
R1297 a_n1236_n9479.n47 a_n1236_n9479.n45 0.459739
R1298 a_n1236_n9479.n49 a_n1236_n9479.n48 0.459739
R1299 a_n1236_n9479.n62 a_n1236_n9479.n37 0.451587
R1300 a_n1236_n9479.n64 a_n1236_n9479.n63 0.451587
R1301 a_n1236_n9479.n54 a_n1236_n9479.n8 0.408833
R1302 a_n1236_n9479.n30 a_n1236_n9479.n28 0.405391
R1303 a_n1236_n9479.n32 a_n1236_n9479.n31 0.405391
R1304 a_n1236_n9479.n73 a_n1236_n9479.n12 0.395292
R1305 a_n1236_n9479.n66 a_n1236_n9479.n10 0.395292
R1306 a_n1236_n9479.n73 a_n1236_n9479.n36 0.143208
R1307 a_n1236_n9479.n68 a_n1236_n9479.n66 0.143208
R1308 2nd_3_OTA_0.vd4.n0 2nd_3_OTA_0.vd4.t11 82.3324
R1309 2nd_3_OTA_0.vd4.n0 2nd_3_OTA_0.vd4.t8 81.6762
R1310 2nd_3_OTA_0.vd4.n0 2nd_3_OTA_0.vd4.t12 81.6762
R1311 2nd_3_OTA_0.vd4.n0 2nd_3_OTA_0.vd4.t10 81.4249
R1312 2nd_3_OTA_0.vd4.n4 2nd_3_OTA_0.vd4.t6 72.7606
R1313 2nd_3_OTA_0.vd4 2nd_3_OTA_0.vd4.t4 71.6732
R1314 2nd_3_OTA_0.vd4 2nd_3_OTA_0.vd4.n5 62.243
R1315 2nd_3_OTA_0.vd4.n1 2nd_3_OTA_0.vd4.t7 19.4751
R1316 2nd_3_OTA_0.vd4.n1 2nd_3_OTA_0.vd4.t1 18.6511
R1317 2nd_3_OTA_0.vd4.n3 2nd_3_OTA_0.vd4.n2 15.6099
R1318 2nd_3_OTA_0.vd4.n5 2nd_3_OTA_0.vd4.t5 11.6005
R1319 2nd_3_OTA_0.vd4.n5 2nd_3_OTA_0.vd4.t3 11.6005
R1320 2nd_3_OTA_0.vd4 2nd_3_OTA_0.vd4.t9 4.23179
R1321 2nd_3_OTA_0.vd4 2nd_3_OTA_0.vd4.n4 2.90758
R1322 2nd_3_OTA_0.vd4 2nd_3_OTA_0.vd4.n0 2.2205
R1323 2nd_3_OTA_0.vd4.n2 2nd_3_OTA_0.vd4.t2 1.90483
R1324 2nd_3_OTA_0.vd4.n2 2nd_3_OTA_0.vd4.t0 1.90483
R1325 2nd_3_OTA_0.vd4.n3 2nd_3_OTA_0.vd4.n1 1.32214
R1326 2nd_3_OTA_0.vd4.n4 2nd_3_OTA_0.vd4.n3 1.28407
R1327 a_7434_1657.n9 a_7434_1657.t12 387.31
R1328 a_7434_1657.n10 a_7434_1657.t5 96.3265
R1329 a_7434_1657.n6 a_7434_1657.t7 96.3265
R1330 a_7434_1657.n3 a_7434_1657.n8 84.9005
R1331 a_7434_1657.n5 a_7434_1657.t10 35.0885
R1332 a_7434_1657.n5 a_7434_1657.t9 34.5018
R1333 a_7434_1657.t4 a_7434_1657.n9 32.649
R1334 a_7434_1657.n7 a_7434_1657.n6 0.971171
R1335 a_7434_1657.n10 a_7434_1657.t4 28.9361
R1336 a_7434_1657.n11 a_7434_1657.n5 28.9216
R1337 a_7434_1657.t0 a_7434_1657.n3 28.1453
R1338 a_7434_1657.n2 a_7434_1657.t2 13.2766
R1339 a_7434_1657.n7 a_7434_1657.t6 13.4238
R1340 a_7434_1657.n8 a_7434_1657.t3 11.4265
R1341 a_7434_1657.n8 a_7434_1657.t1 11.4265
R1342 a_7434_1657.n0 a_7434_1657.n7 7.07514
R1343 a_7434_1657.n1 a_7434_1657.n0 2.67922
R1344 a_7434_1657.n11 a_7434_1657.t8 5.8005
R1345 a_7434_1657.t11 a_7434_1657.n11 5.8005
R1346 a_7434_1657.n1 a_7434_1657.n2 1.64285
R1347 a_7434_1657.n4 a_7434_1657.n6 5.19734
R1348 a_7434_1657.n5 a_7434_1657.n3 3.73846
R1349 a_7434_1657.n9 a_7434_1657.n0 3.7305
R1350 a_7434_1657.n4 a_7434_1657.n10 3.46037
R1351 a_7434_1657.n2 a_7434_1657.n3 1.08359
R1352 a_7434_1657.n5 a_7434_1657.n4 1.8052
R1353 a_7434_1657.n1 a_7434_1657.t0 27.348
R1354 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd2.t2 134.761
R1355 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd2.t3 134.73
R1356 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd2.t5 122.688
R1357 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd2.t8 122.213
R1358 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd2.t6 122.213
R1359 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd2.t7 121.831
R1360 2nd_3_OTA_0.vd2.t4 2nd_3_OTA_0.vd2.t1 26.2097
R1361 2nd_3_OTA_0.vd2.t1 2nd_3_OTA_0.vd2.t0 19.2526
R1362 a_n1050_166.n4 a_n1050_166.t0 36.4777
R1363 a_n1050_166.n5 a_n1050_166.t1 35.4327
R1364 a_n1050_166.n4 a_n1050_166.n3 31.3519
R1365 a_n1050_166.n8 a_n1050_166.n7 18.3035
R1366 a_n1050_166.n2 a_n1050_166.n1 18.303
R1367 a_n1050_166.n9 a_n1050_166.n8 17.2098
R1368 a_n1050_166.n2 a_n1050_166.n0 17.208
R1369 a_n1050_166.n6 a_n1050_166.n2 8.938
R1370 a_n1050_166.n3 a_n1050_166.t3 4.08121
R1371 a_n1050_166.n3 a_n1050_166.t5 4.08121
R1372 a_n1050_166.n8 a_n1050_166.n6 3.05142
R1373 a_n1050_166.n6 a_n1050_166.n5 2.2455
R1374 a_n1050_166.n1 a_n1050_166.t7 1.90483
R1375 a_n1050_166.n1 a_n1050_166.t11 1.90483
R1376 a_n1050_166.n0 a_n1050_166.t4 1.90483
R1377 a_n1050_166.n0 a_n1050_166.t9 1.90483
R1378 a_n1050_166.n7 a_n1050_166.t2 1.90483
R1379 a_n1050_166.n7 a_n1050_166.t8 1.90483
R1380 a_n1050_166.t10 a_n1050_166.n9 1.90483
R1381 a_n1050_166.n9 a_n1050_166.t6 1.90483
R1382 a_n1050_166.n5 a_n1050_166.n4 1.0455
R1383 vcc.n213 vcc.n19 17565.9
R1384 vcc.n215 vcc.n19 17565.9
R1385 vcc.n215 vcc.n20 17562.4
R1386 vcc.n213 vcc.n20 17562.4
R1387 vcc.n8 vcc.n5 16027.1
R1388 vcc.n10 vcc.n5 16027.1
R1389 vcc.n8 vcc.n6 16027.1
R1390 vcc.n10 vcc.n6 16027.1
R1391 vcc.n156 vcc.n57 12420
R1392 vcc.n156 vcc.n46 12420
R1393 vcc.n158 vcc.n57 12416.5
R1394 vcc.n158 vcc.n46 12416.5
R1395 vcc.n204 vcc.n34 6349.41
R1396 vcc.n204 vcc.n35 6349.41
R1397 vcc.n202 vcc.n34 6349.41
R1398 vcc.n202 vcc.n35 6349.41
R1399 vcc.n144 vcc.n56 4698.77
R1400 vcc.n94 vcc.n91 3045.88
R1401 vcc.n97 vcc.n91 3045.88
R1402 vcc.n97 vcc.n92 3045.88
R1403 vcc.n135 vcc.n70 2701.93
R1404 vcc.n131 vcc.n72 2372.5
R1405 vcc.n72 vcc.n71 2327.31
R1406 vcc.n103 vcc.n88 2089.41
R1407 vcc.n106 vcc.n87 2089.41
R1408 vcc.n110 vcc.n79 2089.41
R1409 vcc.n113 vcc.n78 2089.41
R1410 vcc.n120 vcc.n119 2089.41
R1411 vcc.n122 vcc.n75 2089.41
R1412 vcc.n177 vcc.n54 2071.76
R1413 vcc.n171 vcc.n162 2071.76
R1414 vcc.n169 vcc.n55 1443.53
R1415 vcc.n169 vcc.n164 1443.53
R1416 vcc.n10 vcc.t37 1353.8
R1417 vcc.t41 vcc.n8 1317.74
R1418 vcc.n9 vcc.t41 1196.03
R1419 vcc.t37 vcc.n9 1159.97
R1420 vcc.n165 vcc.n164 628.236
R1421 vcc.n164 vcc.n54 628.236
R1422 vcc.n171 vcc.n55 628.236
R1423 vcc.n175 vcc.n55 628.236
R1424 vcc.n66 vcc.n65 599.49
R1425 vcc.n7 vcc.n4 415.628
R1426 vcc.n133 vcc.t23 413.37
R1427 vcc.t7 vcc.t9 412.942
R1428 vcc.t11 vcc.t5 412.942
R1429 vcc.n11 vcc.n4 405.284
R1430 vcc.t23 vcc.t19 387.817
R1431 vcc.t9 vcc.n57 319.411
R1432 vcc.t5 vcc.n46 315.507
R1433 vcc.n104 vcc.n87 290.354
R1434 vcc.n105 vcc.n88 290.354
R1435 vcc.n111 vcc.n78 290.354
R1436 vcc.n112 vcc.n79 290.354
R1437 vcc.n122 vcc.n121 290.354
R1438 vcc.n119 vcc.n118 290.354
R1439 vcc.n128 vcc.n127 285.889
R1440 vcc.n132 vcc.n70 268.555
R1441 vcc.n189 vcc.n188 259.036
R1442 vcc.n130 vcc.n129 253.067
R1443 vcc.n129 vcc.n128 248.246
R1444 vcc.n81 vcc.t31 231.379
R1445 vcc.n142 vcc.t36 231.287
R1446 vcc.n61 vcc.t18 231.287
R1447 vcc.n83 vcc.t22 231.287
R1448 vcc.n82 vcc.t16 231.273
R1449 vcc.t25 vcc.t0 216.05
R1450 vcc.t28 vcc.t2 216.05
R1451 vcc.n212 vcc.n16 209.422
R1452 vcc.n157 vcc.t11 208.423
R1453 vcc.n157 vcc.t7 204.519
R1454 vcc.n141 vcc.n62 202.453
R1455 vcc.n7 vcc.n3 183.016
R1456 vcc.n135 vcc.n134 182.202
R1457 vcc.n97 vcc.t15 178.327
R1458 vcc.n12 vcc.n11 176.572
R1459 vcc.t13 vcc.n170 176.514
R1460 vcc.n170 vcc.t47 176.514
R1461 vcc.t0 vcc.n34 174.992
R1462 vcc.t2 vcc.n35 174.992
R1463 vcc.n95 vcc.n94 174.803
R1464 vcc.n177 vcc.n176 173.517
R1465 vcc.n163 vcc.n162 173.517
R1466 vcc.n72 vcc.t32 172.579
R1467 vcc.n173 vcc.n172 166.4
R1468 vcc.n160 vcc.n159 161.126
R1469 vcc.n217 vcc.n17 157.375
R1470 vcc.n168 vcc.n167 153.976
R1471 vcc.n168 vcc.n52 146.825
R1472 vcc.n98 vcc.n90 128.709
R1473 vcc.n166 vcc.n161 124.802
R1474 vcc.n2 vcc.n0 120.891
R1475 vcc.n2 vcc.n1 119.76
R1476 vcc.n130 vcc.n126 118.385
R1477 vcc.n30 vcc.n29 116.722
R1478 vcc.n216 vcc.n18 115.912
R1479 vcc.n99 vcc.n98 115.841
R1480 vcc.n217 vcc.n216 108.909
R1481 vcc.n203 vcc.t25 108.025
R1482 vcc.n203 vcc.t28 108.025
R1483 vcc.n189 vcc.n47 104.57
R1484 vcc.n117 vcc.n73 101.912
R1485 vcc.n51 vcc.t14 98.0045
R1486 vcc.n51 vcc.t48 97.6911
R1487 vcc.n178 vcc.n53 95.9841
R1488 vcc.n25 vcc.n24 87.9664
R1489 vcc.n25 vcc.n18 87.7954
R1490 vcc.n182 vcc.n50 87.2408
R1491 vcc.n185 vcc.n184 87.2408
R1492 vcc.n44 vcc.n43 87.1446
R1493 vcc.n149 vcc.n60 87.1446
R1494 vcc.n160 vcc.n56 85.5143
R1495 vcc.n117 vcc.n116 82.438
R1496 vcc.n108 vcc.n76 73.7015
R1497 vcc.n115 vcc.n76 72.4513
R1498 vcc.n38 vcc.n37 71.8902
R1499 vcc.t27 vcc.n213 71.3347
R1500 vcc.n201 vcc.n36 70.7824
R1501 vcc.n167 vcc.n166 67.0123
R1502 vcc.n167 vcc.n53 67.0123
R1503 vcc.n172 vcc.n161 65.892
R1504 vcc.n208 vcc.n21 65.6211
R1505 vcc.n107 vcc.n80 64.6513
R1506 vcc.n100 vcc.n80 64.1322
R1507 vcc.n128 vcc.n71 61.6672
R1508 vcc.n172 vcc.n171 61.6672
R1509 vcc.n171 vcc.t13 61.6672
R1510 vcc.n54 vcc.n53 61.6672
R1511 vcc.t47 vcc.n54 61.6672
R1512 vcc.n166 vcc.n165 61.6672
R1513 vcc.n175 vcc.n174 61.6672
R1514 vcc.n215 vcc.t40 60.8049
R1515 vcc.n126 vcc.n125 58.2536
R1516 vcc.n146 vcc.n145 57.394
R1517 vcc.n65 vcc.t33 57.1305
R1518 vcc.n65 vcc.t34 57.1305
R1519 vcc.n134 vcc.n71 56.2313
R1520 vcc.n212 vcc.n211 55.3321
R1521 vcc.n176 vcc.n175 54.8697
R1522 vcc.n165 vcc.n163 54.8697
R1523 vcc.t30 vcc.t27 53.6285
R1524 vcc.t40 vcc.t4 53.6285
R1525 vcc.n205 vcc.n33 50.9389
R1526 vcc.n131 vcc.n130 46.2505
R1527 vcc.n93 vcc.n90 45.8455
R1528 vcc.n133 vcc.t32 43.4751
R1529 vcc.n124 vcc.n73 36.2672
R1530 vcc.n155 vcc.n58 35.1478
R1531 vcc.n132 vcc.n131 33.6572
R1532 vcc.n41 vcc.n39 32.1789
R1533 vcc.t4 vcc.n214 32.0794
R1534 vcc.n41 vcc.n40 32.0774
R1535 vcc.n91 vcc.n90 30.8338
R1536 vcc.n96 vcc.n91 30.8338
R1537 vcc.n103 vcc.n102 30.8338
R1538 vcc.n92 vcc.n89 30.8338
R1539 vcc.n75 vcc.n73 30.8338
R1540 vcc.n126 vcc.n70 30.8338
R1541 vcc.n120 vcc.n74 30.8338
R1542 vcc.n114 vcc.n113 30.8338
R1543 vcc.n110 vcc.n109 30.8338
R1544 vcc.n107 vcc.n106 30.8338
R1545 vcc.n30 vcc.n21 30.7043
R1546 vcc.n206 vcc.n205 30.0503
R1547 vcc.n206 vcc.n32 29.6052
R1548 vcc.t19 vcc.n132 29.2303
R1549 vcc.n95 vcc.n92 28.7736
R1550 vcc.n62 vcc.t20 28.5655
R1551 vcc.n62 vcc.t24 28.5655
R1552 vcc.n104 vcc.n103 26.1635
R1553 vcc.n111 vcc.n110 26.1635
R1554 vcc.n113 vcc.n112 26.1635
R1555 vcc.n121 vcc.n120 26.1635
R1556 vcc.n118 vcc.n75 26.1635
R1557 vcc.n106 vcc.n105 26.1635
R1558 vcc.n146 vcc.n144 24.2792
R1559 vcc.n119 vcc.n117 23.1311
R1560 vcc.n87 vcc.n80 23.1255
R1561 vcc.n101 vcc.n88 23.1255
R1562 vcc.n79 vcc.n76 23.1255
R1563 vcc.n123 vcc.n122 23.1255
R1564 vcc.n78 vcc.n77 23.1255
R1565 vcc.n102 vcc.n101 22.5272
R1566 vcc.n214 vcc.t30 21.5497
R1567 vcc.n162 vcc.n161 18.5005
R1568 vcc.n178 vcc.n177 18.5005
R1569 vcc.n169 vcc.n168 18.5005
R1570 vcc.n170 vcc.n169 18.5005
R1571 vcc.n93 vcc.n89 18.4652
R1572 vcc.n179 vcc.n178 18.1802
R1573 vcc.n179 vcc.n52 17.9947
R1574 vcc.n1 vcc.t42 15.8699
R1575 vcc.n1 vcc.t38 15.8699
R1576 vcc.n0 vcc.t43 15.8699
R1577 vcc.n0 vcc.t39 15.8699
R1578 vcc.n137 vcc.n64 14.6377
R1579 vcc.n127 vcc.n69 14.5701
R1580 vcc.n137 vcc.n136 12.7273
R1581 vcc.n125 vcc.n124 12.0598
R1582 vcc.n159 vcc.n48 11.6663
R1583 vcc.n129 vcc.n72 11.563
R1584 vcc.n50 vcc.t49 11.4265
R1585 vcc.n50 vcc.t8 11.4265
R1586 vcc.n184 vcc.t12 11.4265
R1587 vcc.n184 vcc.t44 11.4265
R1588 vcc.n43 vcc.t46 11.4265
R1589 vcc.n43 vcc.t6 11.4265
R1590 vcc.n60 vcc.t10 11.4265
R1591 vcc.n60 vcc.t45 11.4265
R1592 vcc.n98 vcc.n97 10.8829
R1593 vcc.n94 vcc.n93 10.8829
R1594 vcc.n124 vcc.n123 10.3636
R1595 vcc.n11 vcc.n10 10.2783
R1596 vcc.n8 vcc.n7 10.2783
R1597 vcc.n109 vcc.n77 9.97982
R1598 vcc.n123 vcc.n74 9.86377
R1599 vcc.n116 vcc.n115 9.85683
R1600 vcc.n114 vcc.n77 9.83647
R1601 vcc.n134 vcc.n133 9.79085
R1602 vcc.n100 vcc.n99 9.73877
R1603 vcc.n139 vcc.n64 9.6823
R1604 vcc.n108 vcc.n107 9.62493
R1605 vcc.n101 vcc.n86 9.59483
R1606 vcc.n67 vcc 9.58101
R1607 vcc.n29 vcc.n28 9.34567
R1608 vcc.n59 vcc.n58 9.3005
R1609 vcc.n152 vcc.n47 9.3005
R1610 vcc.n49 vcc.n48 9.3005
R1611 vcc.n200 vcc.n199 9.3005
R1612 vcc.n209 vcc.n208 9.3005
R1613 vcc.n26 vcc.n25 9.3005
R1614 vcc.t15 vcc.n96 8.9954
R1615 vcc.n37 vcc.n35 8.04398
R1616 vcc.n36 vcc.n34 8.04398
R1617 vcc.n136 vcc.n135 7.4005
R1618 vcc vcc.n141 7.20708
R1619 vcc.n202 vcc.n201 7.11588
R1620 vcc.n203 vcc.n202 7.11588
R1621 vcc.n205 vcc.n204 7.11588
R1622 vcc.n204 vcc.n203 7.11588
R1623 vcc.n211 vcc.n21 6.56253
R1624 vcc.n174 vcc.n173 5.75273
R1625 vcc.n190 vcc.n46 5.60656
R1626 vcc.n145 vcc.n57 5.60656
R1627 vcc.n24 vcc.n20 5.44168
R1628 vcc.n214 vcc.n20 5.44168
R1629 vcc.n19 vcc.n17 5.44168
R1630 vcc.n214 vcc.n19 5.44168
R1631 vcc.t13 vcc.n163 5.16575
R1632 vcc.n176 vcc.t47 5.16575
R1633 vcc.n201 vcc.n200 4.82369
R1634 vcc.n173 vcc.n160 4.58844
R1635 vcc.n152 vcc.n151 4.5005
R1636 vcc.n183 vcc.n49 4.5005
R1637 vcc.n36 vcc.n33 4.48345
R1638 vcc.n29 vcc.n22 4.42232
R1639 vcc.n105 vcc.t21 4.28573
R1640 vcc.t21 vcc.n104 4.28573
R1641 vcc.n118 vcc.t35 4.28573
R1642 vcc.n121 vcc.t35 4.28573
R1643 vcc.n112 vcc.t17 4.28573
R1644 vcc.t17 vcc.n111 4.28573
R1645 vcc vcc.n143 4.12557
R1646 vcc.n39 vcc.t1 4.08121
R1647 vcc.n39 vcc.t26 4.08121
R1648 vcc.n40 vcc.t29 4.08121
R1649 vcc.n40 vcc.t3 4.08121
R1650 vcc.n194 vcc.n42 3.98496
R1651 vcc.n187 vcc.n45 3.8313
R1652 vcc.n145 vcc.n56 3.22115
R1653 vcc.n180 vcc.n49 3.09113
R1654 vcc.n159 vcc.n158 2.68166
R1655 vcc.n158 vcc.n157 2.68166
R1656 vcc.n156 vcc.n155 2.68166
R1657 vcc.n157 vcc.n156 2.68166
R1658 vcc.n185 vcc.n42 2.55635
R1659 vcc.n200 vcc.n38 1.94833
R1660 vcc.n28 vcc.n27 1.87667
R1661 vcc.n24 vcc.n22 1.86232
R1662 vcc.n193 vcc.n192 1.85463
R1663 vcc.n219 vcc.n218 1.85361
R1664 vcc.n152 vcc.n45 1.78294
R1665 vcc.n96 vcc.n95 1.7705
R1666 vcc.n182 vcc.n181 1.688
R1667 vcc.n213 vcc.n212 1.66717
R1668 vcc.n216 vcc.n215 1.66717
R1669 vcc.n6 vcc.n4 1.63767
R1670 vcc.n9 vcc.n6 1.63767
R1671 vcc.n5 vcc.n3 1.63767
R1672 vcc.n9 vcc.n5 1.63767
R1673 vcc.n85 vcc.n81 1.62503
R1674 vcc.n207 vcc.n206 1.6211
R1675 vcc.n188 vcc.n48 1.45873
R1676 vcc.n15 vcc.n14 1.41806
R1677 vcc.n183 vcc.n182 1.27935
R1678 vcc.n13 vcc 1.27612
R1679 vcc.n221 vcc.n15 1.21641
R1680 vcc.n17 vcc.n16 1.20392
R1681 vcc.n14 vcc.n2 1.20189
R1682 vcc.n37 vcc.n32 1.19816
R1683 vcc.n147 vcc.n59 1.19668
R1684 vcc.n154 vcc.n47 1.19015
R1685 vcc.n147 vcc.n146 1.11733
R1686 vcc.n144 vcc.n58 1.05462
R1687 vcc.n83 vcc.n82 1.00136
R1688 vcc.n210 vcc.n209 0.985286
R1689 vcc.n26 vcc.n23 0.96321
R1690 vcc.n186 vcc.n185 0.963107
R1691 vcc.n174 vcc.n52 0.933293
R1692 vcc.n198 vcc.n197 0.928261
R1693 vcc.n210 vcc.n30 0.875256
R1694 vcc.n211 vcc.n210 0.862026
R1695 vcc.n195 vcc.n194 0.838031
R1696 vcc.n138 vcc.n68 0.813514
R1697 vcc.n153 vcc.n59 0.780009
R1698 vcc.n27 vcc.n26 0.758322
R1699 vcc.n221 vcc.n220 0.680786
R1700 vcc.n136 vcc.n69 0.649348
R1701 vcc.n148 vcc.n147 0.641762
R1702 vcc.n84 vcc.n83 0.612135
R1703 vcc.n190 vcc.n189 0.603552
R1704 vcc.n85 vcc.n84 0.595437
R1705 vcc.n180 vcc.n179 0.58175
R1706 vcc.n196 vcc.n195 0.539263
R1707 vcc.n143 vcc.n61 0.529588
R1708 vcc.n12 vcc.n3 0.492808
R1709 vcc.n197 vcc.n196 0.445398
R1710 vcc.n193 vcc.n44 0.41511
R1711 vcc.n149 vcc.n148 0.407233
R1712 vcc.n84 vcc.n61 0.403016
R1713 vcc.n220 vcc 0.390072
R1714 vcc.n138 vcc.n137 0.358192
R1715 vcc.n150 vcc.n149 0.347903
R1716 vcc.n27 vcc.n18 0.342518
R1717 vcc.n127 vcc.n68 0.332643
R1718 vcc.n195 vcc.n33 0.321789
R1719 vcc.n82 vcc.n81 0.319213
R1720 vcc.n151 vcc.n44 0.314461
R1721 vcc.n155 vcc.n154 0.2565
R1722 vcc.n181 vcc.n180 0.2505
R1723 vcc.n69 vcc.n63 0.239152
R1724 vcc.n125 vcc.n64 0.237537
R1725 vcc.n99 vcc.n89 0.228778
R1726 vcc.n109 vcc.n108 0.212205
R1727 vcc.n143 vcc.n142 0.180531
R1728 vcc.n140 vcc.n63 0.163235
R1729 vcc.n140 vcc.n139 0.1505
R1730 vcc.n68 vcc.n67 0.1505
R1731 vcc.n191 vcc.n190 0.1505
R1732 vcc.n188 vcc.n187 0.148119
R1733 vcc.n208 vcc.n207 0.137839
R1734 vcc.n181 vcc.n51 0.133423
R1735 vcc.n197 vcc.n32 0.129667
R1736 vcc.n23 vcc.n22 0.129667
R1737 vcc.n13 vcc.n12 0.123496
R1738 vcc.n107 vcc.n86 0.114495
R1739 vcc.n66 vcc.n63 0.111978
R1740 vcc.n198 vcc.n38 0.103833
R1741 vcc.n218 vcc.n217 0.0994362
R1742 vcc vcc.n221 0.0953661
R1743 vcc.n219 vcc.n16 0.0866111
R1744 vcc.n115 vcc.n114 0.0831873
R1745 vcc.n102 vcc.n100 0.0819249
R1746 vcc.n86 vcc.n85 0.0678913
R1747 vcc.n192 vcc.n191 0.0666765
R1748 vcc.n187 vcc.n186 0.0638803
R1749 vcc.n142 vcc 0.0571038
R1750 vcc.n67 vcc.n66 0.0519512
R1751 vcc.n116 vcc.n74 0.0501124
R1752 vcc.n199 vcc.n41 0.047375
R1753 vcc.n148 vcc 0.0443375
R1754 vcc.n218 vcc.n15 0.0429528
R1755 vcc.n220 vcc.n219 0.038
R1756 vcc.n139 vcc.n138 0.037915
R1757 vcc.n194 vcc.n193 0.0364015
R1758 vcc.n207 vcc.n31 0.0341957
R1759 vcc.n141 vcc.n140 0.0303556
R1760 vcc.n154 vcc.n153 0.0274565
R1761 vcc.n153 vcc.n152 0.0266936
R1762 vcc.n151 vcc.n150 0.0261494
R1763 vcc.n192 vcc.n42 0.0233659
R1764 vcc.n199 vcc.n198 0.0216694
R1765 vcc.n187 vcc.n49 0.0211422
R1766 vcc.n196 vcc.n31 0.020648
R1767 vcc.n186 vcc.n183 0.0197308
R1768 vcc.n191 vcc.n45 0.0144018
R1769 vcc.n14 vcc.n13 0.0133125
R1770 vcc.n153 vcc.n150 0.0121883
R1771 vcc.n209 vcc.n31 0.00255592
R1772 vcc.n28 vcc.n23 0.00155302
R1773 vin_p.n0 vin_p.t1 21.6012
R1774 vin_p.n0 vin_p.t0 8.85318
R1775 vin_p vin_p.n0 2.55816
R1776 vo3.n0 vo3.t0 98.4603
R1777 vo3.n0 vo3.t2 88.6727
R1778 vo3.n1 vo3.t1 46.53
R1779 vo3.n1 vo3.n0 0.203972
R1780 vo3 vo3.n1 0.107444
R1781 2nd_3_OTA_0.vb1.n1 2nd_3_OTA_0.vb1.n2 71.7516
R1782 2nd_3_OTA_0.vb1.n1 2nd_3_OTA_0.vb1.n3 70.9453
R1783 2nd_3_OTA_0.vb1.n1 2nd_3_OTA_0.vb1.n4 70.9453
R1784 2nd_3_OTA_0.vb1.n0 2nd_3_OTA_0.vb1.t8 68.1062
R1785 2nd_3_OTA_0.vb1.n0 2nd_3_OTA_0.vb1.t9 67.5138
R1786 2nd_3_OTA_0.vb1.n0 2nd_3_OTA_0.vb1.t7 67.5138
R1787 2nd_3_OTA_0.vb1.n0 2nd_3_OTA_0.vb1.t6 67.5138
R1788 2nd_3_OTA_0.vb1.n2 2nd_3_OTA_0.vb1.t0 17.4005
R1789 2nd_3_OTA_0.vb1.n2 2nd_3_OTA_0.vb1.t2 17.4005
R1790 2nd_3_OTA_0.vb1.n3 2nd_3_OTA_0.vb1.t3 17.4005
R1791 2nd_3_OTA_0.vb1.n3 2nd_3_OTA_0.vb1.t1 17.4005
R1792 2nd_3_OTA_0.vb1.n4 2nd_3_OTA_0.vb1.t4 17.4005
R1793 2nd_3_OTA_0.vb1.n4 2nd_3_OTA_0.vb1.t5 17.4005
R1794 2nd_3_OTA_0.vb1 2nd_3_OTA_0.vb1.n0 10.0205
R1795 2nd_3_OTA_0.vb1 2nd_3_OTA_0.vb1.n1 8.74264
R1796 OTA_vref_0.OTA_vref_stage2_0.vr.n4 OTA_vref_0.OTA_vref_stage2_0.vr.t1 651.943
R1797 OTA_vref_0.OTA_vref_stage2_0.vr.n22 OTA_vref_0.OTA_vref_stage2_0.vr.t3 651.74
R1798 OTA_vref_0.OTA_vref_stage2_0.vr.n24 OTA_vref_0.OTA_vref_stage2_0.vr.t23 60.1752
R1799 OTA_vref_0.OTA_vref_stage2_0.vr.n23 OTA_vref_0.OTA_vref_stage2_0.vr.t22 60.1752
R1800 OTA_vref_0.OTA_vref_stage2_0.vr.n14 OTA_vref_0.OTA_vref_stage2_0.vr.t17 28.5589
R1801 OTA_vref_0.OTA_vref_stage2_0.vr.n18 OTA_vref_0.OTA_vref_stage2_0.vr.t7 27.6016
R1802 OTA_vref_0.OTA_vref_stage2_0.vr.n0 OTA_vref_0.OTA_vref_stage2_0.vr.t25 26.8562
R1803 OTA_vref_0.OTA_vref_stage2_0.vr.n0 OTA_vref_0.OTA_vref_stage2_0.vr.t26 26.0492
R1804 OTA_vref_0.OTA_vref_stage2_0.vr.n1 OTA_vref_0.OTA_vref_stage2_0.vr.t21 26.0492
R1805 OTA_vref_0.OTA_vref_stage2_0.vr.n2 OTA_vref_0.OTA_vref_stage2_0.vr.t24 26.0492
R1806 OTA_vref_0.OTA_vref_stage2_0.vr.n3 OTA_vref_0.OTA_vref_stage2_0.vr.t20 26.0492
R1807 OTA_vref_0.OTA_vref_stage2_0.vr.n9 OTA_vref_0.OTA_vref_stage2_0.vr.n8 24.2089
R1808 OTA_vref_0.OTA_vref_stage2_0.vr.n14 OTA_vref_0.OTA_vref_stage2_0.vr.n13 23.2516
R1809 OTA_vref_0.OTA_vref_stage2_0.vr.n15 OTA_vref_0.OTA_vref_stage2_0.vr.n12 23.2516
R1810 OTA_vref_0.OTA_vref_stage2_0.vr.n9 OTA_vref_0.OTA_vref_stage2_0.vr.n7 23.2516
R1811 OTA_vref_0.OTA_vref_stage2_0.vr.n10 OTA_vref_0.OTA_vref_stage2_0.vr.n6 23.2516
R1812 OTA_vref_0.OTA_vref_stage2_0.vr.n11 OTA_vref_0.OTA_vref_stage2_0.vr.n5 23.2516
R1813 OTA_vref_0.OTA_vref_stage2_0.vr.n17 OTA_vref_0.OTA_vref_stage2_0.vr.n16 23.2516
R1814 OTA_vref_0.OTA_vref_stage2_0.vr.n4 OTA_vref_0.OTA_vref_stage2_0.vr.t0 23
R1815 OTA_vref_0.OTA_vref_stage2_0.vr.n21 OTA_vref_0.OTA_vref_stage2_0.vr.t2 23
R1816 OTA_vref_0.OTA_vref_stage2_0.vr.n13 OTA_vref_0.OTA_vref_stage2_0.vr.t10 4.3505
R1817 OTA_vref_0.OTA_vref_stage2_0.vr.n13 OTA_vref_0.OTA_vref_stage2_0.vr.t4 4.3505
R1818 OTA_vref_0.OTA_vref_stage2_0.vr.n12 OTA_vref_0.OTA_vref_stage2_0.vr.t13 4.3505
R1819 OTA_vref_0.OTA_vref_stage2_0.vr.n12 OTA_vref_0.OTA_vref_stage2_0.vr.t18 4.3505
R1820 OTA_vref_0.OTA_vref_stage2_0.vr.n8 OTA_vref_0.OTA_vref_stage2_0.vr.t9 4.3505
R1821 OTA_vref_0.OTA_vref_stage2_0.vr.n8 OTA_vref_0.OTA_vref_stage2_0.vr.t16 4.3505
R1822 OTA_vref_0.OTA_vref_stage2_0.vr.n7 OTA_vref_0.OTA_vref_stage2_0.vr.t8 4.3505
R1823 OTA_vref_0.OTA_vref_stage2_0.vr.n7 OTA_vref_0.OTA_vref_stage2_0.vr.t12 4.3505
R1824 OTA_vref_0.OTA_vref_stage2_0.vr.n6 OTA_vref_0.OTA_vref_stage2_0.vr.t6 4.3505
R1825 OTA_vref_0.OTA_vref_stage2_0.vr.n6 OTA_vref_0.OTA_vref_stage2_0.vr.t14 4.3505
R1826 OTA_vref_0.OTA_vref_stage2_0.vr.n5 OTA_vref_0.OTA_vref_stage2_0.vr.t5 4.3505
R1827 OTA_vref_0.OTA_vref_stage2_0.vr.n5 OTA_vref_0.OTA_vref_stage2_0.vr.t15 4.3505
R1828 OTA_vref_0.OTA_vref_stage2_0.vr.n16 OTA_vref_0.OTA_vref_stage2_0.vr.t11 4.3505
R1829 OTA_vref_0.OTA_vref_stage2_0.vr.n16 OTA_vref_0.OTA_vref_stage2_0.vr.t19 4.3505
R1830 OTA_vref_0.OTA_vref_stage2_0.vr.n20 OTA_vref_0.OTA_vref_stage2_0.vr.n19 3.89276
R1831 OTA_vref_0.OTA_vref_stage2_0.vr.n1 OTA_vref_0.OTA_vref_stage2_0.vr.n0 2.80213
R1832 OTA_vref_0.OTA_vref_stage2_0.vr.n3 OTA_vref_0.OTA_vref_stage2_0.vr.n2 2.76952
R1833 OTA_vref_0.OTA_vref_stage2_0.vr.n2 OTA_vref_0.OTA_vref_stage2_0.vr.n1 2.72333
R1834 OTA_vref_0.OTA_vref_stage2_0.vr.n19 OTA_vref_0.OTA_vref_stage2_0.vr.n11 1.06728
R1835 OTA_vref_0.OTA_vref_stage2_0.vr.n10 OTA_vref_0.OTA_vref_stage2_0.vr.n9 0.957816
R1836 OTA_vref_0.OTA_vref_stage2_0.vr.n11 OTA_vref_0.OTA_vref_stage2_0.vr.n10 0.957816
R1837 OTA_vref_0.OTA_vref_stage2_0.vr.n15 OTA_vref_0.OTA_vref_stage2_0.vr.n14 0.957816
R1838 OTA_vref_0.OTA_vref_stage2_0.vr.n17 OTA_vref_0.OTA_vref_stage2_0.vr.n15 0.957816
R1839 OTA_vref_0.OTA_vref_stage2_0.vr.n18 OTA_vref_0.OTA_vref_stage2_0.vr.n17 0.957816
R1840 OTA_vref_0.OTA_vref_stage2_0.vr.n23 OTA_vref_0.OTA_vref_stage2_0.vr.n22 0.712457
R1841 OTA_vref_0.OTA_vref_stage2_0.vr OTA_vref_0.OTA_vref_stage2_0.vr.n24 0.660826
R1842 OTA_vref_0.OTA_vref_stage2_0.vr OTA_vref_0.OTA_vref_stage2_0.vr.n3 0.617348
R1843 OTA_vref_0.OTA_vref_stage2_0.vr.n19 OTA_vref_0.OTA_vref_stage2_0.vr.n18 0.577487
R1844 OTA_vref_0.OTA_vref_stage2_0.vr.n24 OTA_vref_0.OTA_vref_stage2_0.vr.n23 0.36463
R1845 OTA_vref_0.OTA_vref_stage2_0.vr.n21 OTA_vref_0.OTA_vref_stage2_0.vr.n20 0.240616
R1846 OTA_vref_0.OTA_vref_stage2_0.vr.n20 OTA_vref_0.OTA_vref_stage2_0.vr.n4 0.216527
R1847 OTA_vref_0.OTA_vref_stage2_0.vr.n22 OTA_vref_0.OTA_vref_stage2_0.vr.n21 0.206939
R1848 a_11275_n2439.t0 a_11275_n2439.t1 50.1091
R1849 2nd_3_OTA_0.vd1.n0 2nd_3_OTA_0.vd1.t0 138.714
R1850 2nd_3_OTA_0.vd1.n1 2nd_3_OTA_0.vd1.t1 136.073
R1851 2nd_3_OTA_0.vd1.n1 2nd_3_OTA_0.vd1.t6 122.216
R1852 2nd_3_OTA_0.vd1.n1 2nd_3_OTA_0.vd1.t4 122.216
R1853 2nd_3_OTA_0.vd1.n1 2nd_3_OTA_0.vd1.t5 121.828
R1854 2nd_3_OTA_0.vd1.n1 2nd_3_OTA_0.vd1.t7 121.828
R1855 2nd_3_OTA_0.vd1.n0 2nd_3_OTA_0.vd1.t2 19.5045
R1856 2nd_3_OTA_0.vd1.n1 2nd_3_OTA_0.vd1.t3 17.559
R1857 2nd_3_OTA_0.vd1.n1 2nd_3_OTA_0.vd1.n0 11.1867
R1858 3rd_3_OTA_0.vd1 2nd_3_OTA_0.vd1.n1 9.24116
R1859 vin_n.n0 vin_n.t1 21.0692
R1860 vin_n.n0 vin_n.t0 8.85313
R1861 vin_n vin_n.n0 2.40005
C0 a_2382_n6868# a_2470_n5378# 1.04e-19
C1 2nd_3_OTA_0.vd4 2nd_3_OTA_0.vd3 9.480929f
C2 vin_n a_n10077_1624# 1.47482f
C3 a_2382_n5578# a_2382_n6868# 0.154516f
C4 vcc a_2470_n5378# 0.034455f
C5 OTA_vref_0.vb 2nd_3_OTA_0.vd4 0.318281f
C6 a_2382_n6868# OTA_vref_0.OTA_vref_stage2_0.vref0 0.010991f
C7 vcc a_2382_n5578# 0.335707f
C8 a_2382_n6868# a_2382_n8158# 0.154705f
C9 a_2382_n6868# 2nd_3_OTA_0.vb1 1.61373f
C10 vcc OTA_vref_0.OTA_vref_stage2_0.vref0 0.030224f
C11 vcc a_2382_n8158# 0.3278f
C12 vcc 2nd_3_OTA_0.vb1 8.322209f
C13 vin_n vcc 0.018448f
C14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2470_n5378# 6.62e-20
C15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2382_n5578# 0.007176f
C16 OTA_vref_0.vb a_2470_n5378# 0.036384f
C17 a_2382_n5578# OTA_vref_0.vb 3.04e-19
C18 2nd_3_OTA_0.vd3 2nd_3_OTA_0.vb1 0.316815f
C19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage2_0.vref0 16.2573f
C20 2nd_3_OTA_0.vd4 a_2382_n4288# 2.1e-20
C21 a_9040_n3397# vcc 0.101608f
C22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2382_n8158# 0.032619f
C23 OTA_vref_0.vb OTA_vref_0.OTA_vref_stage2_0.vref0 4.32e-19
C24 vcc a_n10077_1624# 5.64e-19
C25 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 2nd_3_OTA_0.vb1 6.15e-19
C26 OTA_vref_0.vb 2nd_3_OTA_0.vb1 0.111837f
C27 vin_n OTA_vref_0.vb 0.605449f
C28 a_9040_n3397# 2nd_3_OTA_0.vd3 1.06971f
C29 vcc a_2382_n6868# 0.318981f
C30 a_2382_n4288# a_2470_n5378# 0.10061f
C31 a_2382_n5578# a_2382_n4288# 0.154422f
C32 a_9040_n3397# OTA_vref_0.vb 0.541253f
C33 a_n10077_1624# OTA_vref_0.vb 0.443825f
C34 a_11847_n1701# vo3 0.159655f
C35 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2382_n6868# 0.009524f
C36 vcc 2nd_3_OTA_0.vd3 4.62835f
C37 a_2470_n7958# OTA_vref_0.OTA_vref_stage2_0.vref0 0.037994f
C38 a_2470_n7958# a_2382_n8158# 1.53765f
C39 a_2470_n7958# 2nd_3_OTA_0.vb1 0.056235f
C40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter vcc 0.512021f
C41 a_11847_n1701# 2nd_3_OTA_0.vd4 1.15e-20
C42 vcc OTA_vref_0.vb 0.434712f
C43 a_2470_n5378# OTA_vref_0.OTA_vref_stage2_0.vr 0.008037f
C44 OTA_vref_0.vb 2nd_3_OTA_0.vd3 0.494477f
C45 a_2382_n5578# OTA_vref_0.OTA_vref_stage2_0.vr 0.334808f
C46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.vb 0.006315f
C47 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vr 2.20674f
C48 a_2382_n8158# OTA_vref_0.OTA_vref_stage2_0.vr 0.33605f
C49 2nd_3_OTA_0.vb1 OTA_vref_0.OTA_vref_stage2_0.vr 0.062593f
C50 vcc a_2382_n4288# 0.368035f
C51 a_2382_n6868# a_2470_n7958# 0.097592f
C52 vcc a_2470_n7958# 0.034292f
C53 2nd_3_OTA_0.vd3 a_2382_n4288# 0.00236f
C54 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2382_n4288# 0.002329f
C55 a_9040_n3397# a_11847_n1701# 0.016974f
C56 OTA_vref_0.vb a_2382_n4288# 1.67298f
C57 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2470_n7958# 0.003419f
C58 vin_p vin_n 2.36446f
C59 a_2382_n6868# OTA_vref_0.OTA_vref_stage2_0.vr 0.341152f
C60 vcc OTA_vref_0.OTA_vref_stage2_0.vr 11.398701f
C61 vin_p a_n10077_1624# 1.68092f
C62 a_11847_n1701# vcc 0.836592f
C63 2nd_3_OTA_0.vd3 OTA_vref_0.OTA_vref_stage2_0.vr 0.001587f
C64 2nd_3_OTA_0.vd4 2nd_3_OTA_0.vb1 0.226739f
C65 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage2_0.vr 9.256969f
C66 a_11847_n1701# 2nd_3_OTA_0.vd3 6.67e-20
C67 OTA_vref_0.vb OTA_vref_0.OTA_vref_stage2_0.vr 0.233485f
C68 a_9040_n3397# vo3 0.004168f
C69 a_2382_n5578# a_2470_n5378# 1.53005f
C70 vin_p vcc 0.018752f
C71 a_2470_n5378# OTA_vref_0.OTA_vref_stage2_0.vref0 0.00151f
C72 a_9040_n3397# 2nd_3_OTA_0.vd4 1.05152f
C73 a_2382_n5578# OTA_vref_0.OTA_vref_stage2_0.vref0 0.011315f
C74 2nd_3_OTA_0.vb1 a_2470_n5378# 0.038035f
C75 a_2382_n5578# 2nd_3_OTA_0.vb1 0.106848f
C76 a_2382_n8158# OTA_vref_0.OTA_vref_stage2_0.vref0 0.112341f
C77 2nd_3_OTA_0.vb1 OTA_vref_0.OTA_vref_stage2_0.vref0 0.006422f
C78 a_2382_n4288# OTA_vref_0.OTA_vref_stage2_0.vr 0.368863f
C79 a_2382_n8158# 2nd_3_OTA_0.vb1 0.034229f
C80 vin_p OTA_vref_0.vb 0.39332f
C81 vo3 vcc 0.594996f
C82 vcc 2nd_3_OTA_0.vd4 4.40467f
C83 a_2470_n7958# OTA_vref_0.OTA_vref_stage2_0.vr 0.008049f
C84 vo3 vss 2.83219f
C85 vin_n vss 15.210062f
C86 vin_p vss 14.908583f
C87 vcc vss 0.224583p
C88 a_2382_n8158# vss 3.83372f
C89 a_2470_n7958# vss 0.471548f
C90 a_2382_n6868# vss 3.70817f
C91 a_2382_n5578# vss 3.70757f
C92 a_2470_n5378# vss 0.471213f
C93 a_2382_n4288# vss 3.74312f
C94 OTA_vref_0.OTA_vref_stage2_0.vref0 vss 14.810505f
C95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter vss 25.278364f
C96 OTA_vref_0.OTA_vref_stage2_0.vr vss 12.014772f
C97 a_11847_n1701# vss 1.4749f
C98 a_9040_n3397# vss 5.75308f
C99 2nd_3_OTA_0.vb1 vss 8.843204f
C100 2nd_3_OTA_0.vd3 vss 48.63614f
C101 2nd_3_OTA_0.vd4 vss 20.133524f
C102 OTA_vref_0.vb vss 17.2421f
C103 a_n10077_1624# vss 3.49104f
C104 vin_n.t1 vss 0.869123f
C105 vin_n.t0 vss 0.457268f
C106 vin_n.n0 vss 1.00705f
C107 2nd_3_OTA_0.vd1.n0 vss 1.9415f
C108 2nd_3_OTA_0.vd1.n1 vss 19.1674f
C109 3rd_3_OTA_0.vd1 vss 37.252304f
C110 2nd_3_OTA_0.vd1.t1 vss 0.043314f
C111 2nd_3_OTA_0.vd1.t0 vss 0.047902f
C112 2nd_3_OTA_0.vd1.t2 vss 0.356063f
C113 2nd_3_OTA_0.vd1.t3 vss 0.217646f
C114 2nd_3_OTA_0.vd1.t5 vss 1.58819f
C115 2nd_3_OTA_0.vd1.t6 vss 1.59871f
C116 2nd_3_OTA_0.vd1.t4 vss 1.59871f
C117 2nd_3_OTA_0.vd1.t7 vss 1.58819f
C118 a_11275_n2439.t1 vss 26.271801f
C119 a_11275_n2439.t0 vss 0.028206f
C120 OTA_vref_0.OTA_vref_stage2_0.vr.t25 vss 0.60782f
C121 OTA_vref_0.OTA_vref_stage2_0.vr.t26 vss 0.584499f
C122 OTA_vref_0.OTA_vref_stage2_0.vr.n0 vss 1.65263f
C123 OTA_vref_0.OTA_vref_stage2_0.vr.t21 vss 0.584499f
C124 OTA_vref_0.OTA_vref_stage2_0.vr.n1 vss 0.976322f
C125 OTA_vref_0.OTA_vref_stage2_0.vr.t24 vss 0.584499f
C126 OTA_vref_0.OTA_vref_stage2_0.vr.n2 vss 0.97502f
C127 OTA_vref_0.OTA_vref_stage2_0.vr.t20 vss 0.584499f
C128 OTA_vref_0.OTA_vref_stage2_0.vr.n3 vss 0.890892f
C129 OTA_vref_0.OTA_vref_stage2_0.vr.t23 vss 0.303436f
C130 OTA_vref_0.OTA_vref_stage2_0.vr.t22 vss 0.303436f
C131 OTA_vref_0.OTA_vref_stage2_0.vr.t3 vss 0.025841f
C132 OTA_vref_0.OTA_vref_stage2_0.vr.t2 vss 0.458739f
C133 OTA_vref_0.OTA_vref_stage2_0.vr.t0 vss 0.458739f
C134 OTA_vref_0.OTA_vref_stage2_0.vr.t1 vss 0.02587f
C135 OTA_vref_0.OTA_vref_stage2_0.vr.n4 vss 0.832695f
C136 OTA_vref_0.OTA_vref_stage2_0.vr.t5 vss 0.054748f
C137 OTA_vref_0.OTA_vref_stage2_0.vr.t15 vss 0.054748f
C138 OTA_vref_0.OTA_vref_stage2_0.vr.n5 vss 0.20797f
C139 OTA_vref_0.OTA_vref_stage2_0.vr.t6 vss 0.054748f
C140 OTA_vref_0.OTA_vref_stage2_0.vr.t14 vss 0.054748f
C141 OTA_vref_0.OTA_vref_stage2_0.vr.n6 vss 0.20797f
C142 OTA_vref_0.OTA_vref_stage2_0.vr.t8 vss 0.054748f
C143 OTA_vref_0.OTA_vref_stage2_0.vr.t12 vss 0.054748f
C144 OTA_vref_0.OTA_vref_stage2_0.vr.n7 vss 0.20797f
C145 OTA_vref_0.OTA_vref_stage2_0.vr.t9 vss 0.054748f
C146 OTA_vref_0.OTA_vref_stage2_0.vr.t16 vss 0.054748f
C147 OTA_vref_0.OTA_vref_stage2_0.vr.n8 vss 0.236203f
C148 OTA_vref_0.OTA_vref_stage2_0.vr.n9 vss 1.66546f
C149 OTA_vref_0.OTA_vref_stage2_0.vr.n10 vss 0.97974f
C150 OTA_vref_0.OTA_vref_stage2_0.vr.n11 vss 1.0171f
C151 OTA_vref_0.OTA_vref_stage2_0.vr.t7 vss 0.276061f
C152 OTA_vref_0.OTA_vref_stage2_0.vr.t13 vss 0.054748f
C153 OTA_vref_0.OTA_vref_stage2_0.vr.t18 vss 0.054748f
C154 OTA_vref_0.OTA_vref_stage2_0.vr.n12 vss 0.20797f
C155 OTA_vref_0.OTA_vref_stage2_0.vr.t10 vss 0.054748f
C156 OTA_vref_0.OTA_vref_stage2_0.vr.t4 vss 0.054748f
C157 OTA_vref_0.OTA_vref_stage2_0.vr.n13 vss 0.20797f
C158 OTA_vref_0.OTA_vref_stage2_0.vr.t17 vss 0.301381f
C159 OTA_vref_0.OTA_vref_stage2_0.vr.n14 vss 1.70977f
C160 OTA_vref_0.OTA_vref_stage2_0.vr.n15 vss 0.97974f
C161 OTA_vref_0.OTA_vref_stage2_0.vr.t11 vss 0.054748f
C162 OTA_vref_0.OTA_vref_stage2_0.vr.t19 vss 0.054748f
C163 OTA_vref_0.OTA_vref_stage2_0.vr.n16 vss 0.20797f
C164 OTA_vref_0.OTA_vref_stage2_0.vr.n17 vss 0.97974f
C165 OTA_vref_0.OTA_vref_stage2_0.vr.n18 vss 0.920416f
C166 OTA_vref_0.OTA_vref_stage2_0.vr.n19 vss 1.68401f
C167 OTA_vref_0.OTA_vref_stage2_0.vr.n20 vss 0.843703f
C168 OTA_vref_0.OTA_vref_stage2_0.vr.n21 vss 0.768139f
C169 OTA_vref_0.OTA_vref_stage2_0.vr.n22 vss 0.122166f
C170 OTA_vref_0.OTA_vref_stage2_0.vr.n23 vss 0.367868f
C171 OTA_vref_0.OTA_vref_stage2_0.vr.n24 vss 0.365806f
C172 2nd_3_OTA_0.vb1.n0 vss 5.75346f
C173 2nd_3_OTA_0.vb1.n1 vss 0.352136f
C174 2nd_3_OTA_0.vb1.t8 vss 0.858318f
C175 2nd_3_OTA_0.vb1.t9 vss 0.846486f
C176 2nd_3_OTA_0.vb1.t7 vss 0.846486f
C177 2nd_3_OTA_0.vb1.t6 vss 0.846486f
C178 2nd_3_OTA_0.vb1.t0 vss 0.007035f
C179 2nd_3_OTA_0.vb1.t2 vss 0.007035f
C180 2nd_3_OTA_0.vb1.n2 vss 0.018857f
C181 2nd_3_OTA_0.vb1.t3 vss 0.007035f
C182 2nd_3_OTA_0.vb1.t1 vss 0.007035f
C183 2nd_3_OTA_0.vb1.n3 vss 0.017824f
C184 2nd_3_OTA_0.vb1.t4 vss 0.007035f
C185 2nd_3_OTA_0.vb1.t5 vss 0.007035f
C186 2nd_3_OTA_0.vb1.n4 vss 0.017824f
C187 vin_p.t1 vss 0.872831f
C188 vin_p.t0 vss 0.458725f
C189 vin_p.n0 vss 1.00306f
C190 vcc.t43 vss 0.004075f
C191 vcc.t39 vss 0.004075f
C192 vcc.n0 vss 0.008942f
C193 vcc.t42 vss 0.004075f
C194 vcc.t38 vss 0.004075f
C195 vcc.n1 vss 0.008515f
C196 vcc.n2 vss 0.094492f
C197 vcc.n3 vss 0.63185f
C198 vcc.n4 vss 0.453088f
C199 vcc.n5 vss 0.120661f
C200 vcc.n6 vss 0.120661f
C201 vcc.n7 vss 0.831817f
C202 vcc.n8 vss 1.4329f
C203 vcc.t41 vss 2.24823f
C204 vcc.n9 vss 2.10607f
C205 vcc.t37 vss 2.24793f
C206 vcc.n10 vss 1.43089f
C207 vcc.n11 vss 0.896155f
C208 vcc.n12 vss 0.800752f
C209 vcc.n13 vss 1.07553f
C210 vcc.n14 vss 0.725808f
C211 vcc.n15 vss 0.660326f
C212 vcc.n16 vss 0.418747f
C213 vcc.n17 vss 0.277315f
C214 vcc.n18 vss 0.741112f
C215 vcc.n19 vss 0.132791f
C216 vcc.n20 vss 0.132765f
C217 vcc.n21 vss 0.605507f
C218 vcc.n22 vss 0.005216f
C219 vcc.n23 vss 0.07734f
C220 vcc.n24 vss 0.075575f
C221 vcc.n25 vss 0.241418f
C222 vcc.n26 vss 0.189413f
C223 vcc.n27 vss 0.285392f
C224 vcc.n28 vss 0.47441f
C225 vcc.n29 vss 0.143663f
C226 vcc.n30 vss 0.478074f
C227 vcc.n31 vss 0.006408f
C228 vcc.n32 vss 0.109866f
C229 vcc.n33 vss 0.855462f
C230 vcc.n34 vss 0.34186f
C231 vcc.n35 vss 0.34186f
C232 vcc.t0 vss 0.545767f
C233 vcc.t25 vss 0.449832f
C234 vcc.n36 vss 0.372515f
C235 vcc.n37 vss 0.25669f
C236 vcc.n38 vss 0.212142f
C237 vcc.t1 vss 0.015848f
C238 vcc.t26 vss 0.015848f
C239 vcc.n39 vss 0.041165f
C240 vcc.t29 vss 0.015848f
C241 vcc.t3 vss 0.015848f
C242 vcc.n40 vss 0.040406f
C243 vcc.n41 vss 0.646562f
C244 vcc.n42 vss 0.127804f
C245 vcc.t46 vss 0.00566f
C246 vcc.t6 vss 0.00566f
C247 vcc.n43 vss 0.012266f
C248 vcc.n44 vss 0.382634f
C249 vcc.n45 vss 0.365143f
C250 vcc.n46 vss 0.963739f
C251 vcc.n47 vss 1.45885f
C252 vcc.n48 vss 0.009991f
C253 vcc.n49 vss 0.1179f
C254 vcc.t49 vss 0.00566f
C255 vcc.t8 vss 0.00566f
C256 vcc.n50 vss 0.012316f
C257 vcc.t14 vss 0.022563f
C258 vcc.t48 vss 0.022382f
C259 vcc.n51 vss 0.118299f
C260 vcc.n52 vss 0.022568f
C261 vcc.n53 vss 0.016393f
C262 vcc.n54 vss 0.010467f
C263 vcc.t47 vss 0.143197f
C264 vcc.n55 vss 0.010153f
C265 vcc.n56 vss 0.069181f
C266 vcc.n57 vss 0.943396f
C267 vcc.t9 vss 1.78421f
C268 vcc.t7 vss 1.50302f
C269 vcc.t5 vss 1.77527f
C270 vcc.t11 vss 1.51252f
C271 vcc.n58 vss 0.79761f
C272 vcc.n59 vss 0.388354f
C273 vcc.t10 vss 0.00566f
C274 vcc.t45 vss 0.00566f
C275 vcc.n60 vss 0.012266f
C276 vcc.t18 vss 0.008487f
C277 vcc.n61 vss 0.099777f
C278 vcc.t36 vss 0.008487f
C279 vcc.t20 vss 0.002264f
C280 vcc.t24 vss 0.002264f
C281 vcc.n62 vss 0.004829f
C282 vcc.n63 vss 0.297858f
C283 vcc.n64 vss 0.085621f
C284 vcc.t33 vss 0.001132f
C285 vcc.t34 vss 0.001132f
C286 vcc.n65 vss 0.002372f
C287 vcc.n66 vss 0.092849f
C288 vcc.n67 vss 0.167974f
C289 vcc.n68 vss 0.110267f
C290 vcc.n69 vss 0.163502f
C291 vcc.n70 vss 0.111054f
C292 vcc.n71 vss 0.044157f
C293 vcc.t32 vss 0.127015f
C294 vcc.n72 vss 0.175771f
C295 vcc.n73 vss 0.025356f
C296 vcc.n74 vss 0.069745f
C297 vcc.n75 vss 0.01621f
C298 vcc.t35 vss 0.180009f
C299 vcc.n76 vss 0.027447f
C300 vcc.n77 vss 0.109405f
C301 vcc.n78 vss 0.123349f
C302 vcc.n79 vss 0.123349f
C303 vcc.n80 vss 0.029346f
C304 vcc.t31 vss 0.008535f
C305 vcc.n81 vss 0.321749f
C306 vcc.t22 vss 0.008487f
C307 vcc.t16 vss 0.008487f
C308 vcc.n82 vss 0.138208f
C309 vcc.n83 vss 0.153912f
C310 vcc.n84 vss 0.319276f
C311 vcc.n85 vss 0.176914f
C312 vcc.n86 vss 0.071269f
C313 vcc.n87 vss 0.123349f
C314 vcc.n88 vss 0.123349f
C315 vcc.n89 vss 0.11909f
C316 vcc.n90 vss 0.099036f
C317 vcc.n91 vss 0.023542f
C318 vcc.n92 vss 0.023542f
C319 vcc.n93 vss 0.283282f
C320 vcc.n94 vss 0.216509f
C321 vcc.n96 vss 0.155553f
C322 vcc.t15 vss 0.148566f
C323 vcc.n97 vss 0.206347f
C324 vcc.n98 vss 0.049103f
C325 vcc.n99 vss 0.21184f
C326 vcc.n100 vss 0.202897f
C327 vcc.n101 vss 0.132849f
C328 vcc.n102 vss 0.047564f
C329 vcc.n103 vss 0.01621f
C330 vcc.t21 vss 0.180009f
C331 vcc.n106 vss 0.01621f
C332 vcc.n107 vss 0.20048f
C333 vcc.n108 vss 0.200676f
C334 vcc.n109 vss 0.070185f
C335 vcc.n110 vss 0.01621f
C336 vcc.t17 vss 0.180009f
C337 vcc.n113 vss 0.01621f
C338 vcc.n114 vss 0.070991f
C339 vcc.n115 vss 0.197547f
C340 vcc.n116 vss 0.195941f
C341 vcc.n117 vss 0.028712f
C342 vcc.n119 vss 0.123351f
C343 vcc.n120 vss 0.01621f
C344 vcc.n122 vss 0.123349f
C345 vcc.n123 vss 0.111372f
C346 vcc.n124 vss 0.132628f
C347 vcc.n125 vss 0.074244f
C348 vcc.n126 vss 0.013276f
C349 vcc.n127 vss 0.264722f
C350 vcc.n128 vss 0.03185f
C351 vcc.n129 vss 0.035677f
C352 vcc.n130 vss 0.026705f
C353 vcc.n131 vss 0.026705f
C354 vcc.n132 vss 0.040493f
C355 vcc.t19 vss 0.091731f
C356 vcc.t23 vss 0.131487f
C357 vcc.n133 vss 0.144827f
C358 vcc.n134 vss 0.068944f
C359 vcc.n135 vss 0.215965f
C360 vcc.n136 vss 0.076568f
C361 vcc.n137 vss 0.155259f
C362 vcc.n138 vss 0.05679f
C363 vcc.n139 vss 0.059208f
C364 vcc.n140 vss 0.087299f
C365 vcc.n141 vss 0.15628f
C366 vcc.n142 vss 0.044913f
C367 vcc.n143 vss 4.31446f
C368 vcc.n144 vss 0.094224f
C369 vcc.n145 vss 0.044408f
C370 vcc.n146 vss 0.084833f
C371 vcc.n147 vss 0.077878f
C372 vcc.n148 vss 0.277515f
C373 vcc.n149 vss 0.394097f
C374 vcc.n150 vss 0.17267f
C375 vcc.n151 vss 0.157191f
C376 vcc.n152 vss 0.596123f
C377 vcc.n153 vss 0.357589f
C378 vcc.n154 vss 0.031851f
C379 vcc.n155 vss 0.780025f
C380 vcc.n156 vss 0.093695f
C381 vcc.n157 vss 1.00518f
C382 vcc.n158 vss 0.093668f
C383 vcc.n159 vss 0.131599f
C384 vcc.n160 vss 0.248041f
C385 vcc.n161 vss 0.040093f
C386 vcc.n162 vss 0.111979f
C387 vcc.n164 vss 0.010153f
C388 vcc.n165 vss 0.010467f
C389 vcc.n166 vss 0.013695f
C390 vcc.n167 vss 0.010153f
C391 vcc.n168 vss 0.010604f
C392 vcc.n169 vss 0.010856f
C393 vcc.n170 vss 0.133123f
C394 vcc.t13 vss 0.143197f
C395 vcc.n171 vss 0.010467f
C396 vcc.n172 vss 0.14043f
C397 vcc.n173 vss 0.07973f
C398 vcc.n174 vss 0.049749f
C399 vcc.n175 vss 0.010467f
C400 vcc.n177 vss 0.111979f
C401 vcc.n178 vss 0.050712f
C402 vcc.n179 vss 0.021008f
C403 vcc.n180 vss 0.186127f
C404 vcc.n181 vss 0.039f
C405 vcc.n182 vss 0.173142f
C406 vcc.n183 vss 0.055488f
C407 vcc.t12 vss 0.00566f
C408 vcc.t44 vss 0.00566f
C409 vcc.n184 vss 0.012316f
C410 vcc.n185 vss 0.199256f
C411 vcc.n186 vss 0.04197f
C412 vcc.n187 vss 0.143462f
C413 vcc.n188 vss 0.204749f
C414 vcc.n189 vss 0.557533f
C415 vcc.n190 vss 0.071534f
C416 vcc.n191 vss 0.046643f
C417 vcc.n192 vss 0.039912f
C418 vcc.n193 vss 0.246993f
C419 vcc.n194 vss 0.48994f
C420 vcc.n195 vss 1.3092f
C421 vcc.n196 vss 0.692498f
C422 vcc.n197 vss 0.270345f
C423 vcc.n198 vss 0.192223f
C424 vcc.n199 vss 0.20619f
C425 vcc.n200 vss 0.015729f
C426 vcc.n201 vss 0.232556f
C427 vcc.n202 vss 0.048176f
C428 vcc.t2 vss 0.545767f
C429 vcc.t28 vss 0.449832f
C430 vcc.n203 vss 0.299888f
C431 vcc.n204 vss 0.048176f
C432 vcc.n205 vss 0.560233f
C433 vcc.n206 vss 0.31532f
C434 vcc.n207 vss 0.011641f
C435 vcc.n208 vss 0.435459f
C436 vcc.n209 vss 0.284788f
C437 vcc.n210 vss 0.436958f
C438 vcc.n211 vss 0.199f
C439 vcc.n212 vss 0.601672f
C440 vcc.n213 vss 2.62577f
C441 vcc.t27 vss 3.10946f
C442 vcc.t30 vss 1.85956f
C443 vcc.n214 vss 1.32653f
C444 vcc.t4 vss 2.12002f
C445 vcc.t40 vss 2.84771f
C446 vcc.n215 vss 2.20306f
C447 vcc.n216 vss 0.3754f
C448 vcc.n217 vss 0.453483f
C449 vcc.n218 vss 0.458572f
C450 vcc.n219 vss 0.47018f
C451 vcc.n220 vss 0.767146f
C452 vcc.n221 vss 0.223998f
C453 a_n1050_166.t6 vss 0.216942f
C454 a_n1050_166.t4 vss 0.216942f
C455 a_n1050_166.t9 vss 0.216942f
C456 a_n1050_166.n0 vss 0.671366f
C457 a_n1050_166.t7 vss 0.216942f
C458 a_n1050_166.t11 vss 0.216942f
C459 a_n1050_166.n1 vss 0.762068f
C460 a_n1050_166.n2 vss 4.7253f
C461 a_n1050_166.t1 vss 0.399519f
C462 a_n1050_166.t3 vss 0.10124f
C463 a_n1050_166.t5 vss 0.10124f
C464 a_n1050_166.n3 vss 0.235864f
C465 a_n1050_166.t0 vss 0.427351f
C466 a_n1050_166.n4 vss 2.07187f
C467 a_n1050_166.n5 vss 1.4064f
C468 a_n1050_166.n6 vss 2.8881f
C469 a_n1050_166.t2 vss 0.216942f
C470 a_n1050_166.t8 vss 0.216942f
C471 a_n1050_166.n7 vss 0.76209f
C472 a_n1050_166.n8 vss 3.54056f
C473 a_n1050_166.n9 vss 0.671495f
C474 a_n1050_166.t10 vss 0.216942f
C475 2nd_3_OTA_0.vd2.t1 vss 38.337997f
C476 2nd_3_OTA_0.vd2.t5 vss 1.328f
C477 2nd_3_OTA_0.vd2.t6 vss 1.32133f
C478 2nd_3_OTA_0.vd2.t8 vss 1.32133f
C479 2nd_3_OTA_0.vd2.t7 vss 1.31275f
C480 2nd_3_OTA_0.vd2.t0 vss 0.353982f
C481 2nd_3_OTA_0.vd2.t2 vss 0.033752f
C482 2nd_3_OTA_0.vd2.t4 vss 0.257087f
C483 2nd_3_OTA_0.vd2.t3 vss 0.03374f
C484 a_7434_1657.n0 vss 1.17962f
C485 a_7434_1657.n1 vss 1.22804f
C486 a_7434_1657.n2 vss 0.281253f
C487 a_7434_1657.t2 vss 1.50909f
C488 a_7434_1657.n3 vss 1.29217f
C489 a_7434_1657.n4 vss 1.58696f
C490 a_7434_1657.n5 vss 3.86795f
C491 a_7434_1657.n6 vss 1.02899f
C492 a_7434_1657.n7 vss 0.64178f
C493 a_7434_1657.t8 vss 0.026714f
C494 a_7434_1657.t12 vss 0.12612f
C495 a_7434_1657.t7 vss 0.081856f
C496 a_7434_1657.t6 vss 1.51857f
C497 a_7434_1657.t3 vss 0.022262f
C498 a_7434_1657.t1 vss 0.022262f
C499 a_7434_1657.n8 vss 0.045353f
C500 a_7434_1657.t0 vss 1.52061f
C501 a_7434_1657.n9 vss 1.63593f
C502 a_7434_1657.t4 vss 1.63702f
C503 a_7434_1657.t5 vss 0.081856f
C504 a_7434_1657.n10 vss 0.711803f
C505 a_7434_1657.t10 vss 0.129672f
C506 a_7434_1657.t9 vss 0.118908f
C507 a_7434_1657.n11 vss 0.078485f
C508 a_7434_1657.t11 vss 0.026714f
C509 2nd_3_OTA_0.vd4.n0 vss 1.19791f
C510 2nd_3_OTA_0.vd4.t11 vss 0.557947f
C511 2nd_3_OTA_0.vd4.t12 vss 0.559799f
C512 2nd_3_OTA_0.vd4.t8 vss 0.559799f
C513 2nd_3_OTA_0.vd4.t10 vss 0.555128f
C514 2nd_3_OTA_0.vd4.t9 vss 16.543098f
C515 2nd_3_OTA_0.vd4.t6 vss 0.04967f
C516 2nd_3_OTA_0.vd4.t1 vss 0.43452f
C517 2nd_3_OTA_0.vd4.t7 vss 0.482932f
C518 2nd_3_OTA_0.vd4.n1 vss 2.53677f
C519 2nd_3_OTA_0.vd4.t2 vss 0.091357f
C520 2nd_3_OTA_0.vd4.t0 vss 0.091357f
C521 2nd_3_OTA_0.vd4.n2 vss 0.253746f
C522 2nd_3_OTA_0.vd4.n3 vss 1.47312f
C523 2nd_3_OTA_0.vd4.n4 vss 1.4592f
C524 2nd_3_OTA_0.vd4.t4 vss 0.044809f
C525 2nd_3_OTA_0.vd4.t5 vss 0.009136f
C526 2nd_3_OTA_0.vd4.t3 vss 0.009136f
C527 2nd_3_OTA_0.vd4.n5 vss 0.054041f
C528 a_n1236_n9479.n0 vss 0.297823f
C529 a_n1236_n9479.n1 vss 0.297439f
C530 a_n1236_n9479.n2 vss 0.29823f
C531 a_n1236_n9479.n3 vss 0.29615f
C532 a_n1236_n9479.n4 vss 0.295296f
C533 a_n1236_n9479.n5 vss 0.585351f
C534 a_n1236_n9479.n6 vss 0.294839f
C535 a_n1236_n9479.n7 vss 0.126637f
C536 a_n1236_n9479.n8 vss 0.297117f
C537 a_n1236_n9479.n9 vss 0.755844f
C538 a_n1236_n9479.n10 vss 0.293675f
C539 a_n1236_n9479.n11 vss 0.295194f
C540 a_n1236_n9479.n12 vss 0.292701f
C541 a_n1236_n9479.n13 vss 0.232375f
C542 a_n1236_n9479.t46 vss 0.036678f
C543 a_n1236_n9479.n14 vss 0.160547f
C544 a_n1236_n9479.n15 vss 0.15275f
C545 a_n1236_n9479.t6 vss 0.428407f
C546 a_n1236_n9479.n16 vss 0.188243f
C547 a_n1236_n9479.t37 vss 0.036678f
C548 a_n1236_n9479.t17 vss 0.036678f
C549 a_n1236_n9479.n17 vss 0.078298f
C550 a_n1236_n9479.n18 vss 0.188647f
C551 a_n1236_n9479.t16 vss 0.428407f
C552 a_n1236_n9479.n19 vss 0.126601f
C553 a_n1236_n9479.t30 vss 0.428407f
C554 a_n1236_n9479.n20 vss 0.191708f
C555 a_n1236_n9479.n21 vss 0.191714f
C556 a_n1236_n9479.n22 vss 0.126636f
C557 a_n1236_n9479.n23 vss 0.252394f
C558 a_n1236_n9479.n24 vss 0.235053f
C559 a_n1236_n9479.t14 vss 0.429053f
C560 a_n1236_n9479.n25 vss 0.501918f
C561 a_n1236_n9479.t15 vss 0.036678f
C562 a_n1236_n9479.t36 vss 0.036678f
C563 a_n1236_n9479.n26 vss 0.078351f
C564 a_n1236_n9479.t39 vss 0.036678f
C565 a_n1236_n9479.t3 vss 0.036678f
C566 a_n1236_n9479.n27 vss 0.078351f
C567 a_n1236_n9479.n28 vss 0.209863f
C568 a_n1236_n9479.n29 vss 0.152512f
C569 a_n1236_n9479.n30 vss 0.210635f
C570 a_n1236_n9479.t2 vss 0.428407f
C571 a_n1236_n9479.n31 vss 0.244957f
C572 a_n1236_n9479.t28 vss 0.428407f
C573 a_n1236_n9479.n32 vss 0.198133f
C574 a_n1236_n9479.n33 vss 0.152497f
C575 a_n1236_n9479.t29 vss 0.036678f
C576 a_n1236_n9479.t45 vss 0.036678f
C577 a_n1236_n9479.n34 vss 0.078351f
C578 a_n1236_n9479.t40 vss 0.036678f
C579 a_n1236_n9479.t7 vss 0.036678f
C580 a_n1236_n9479.n35 vss 0.078353f
C581 a_n1236_n9479.n36 vss 0.224428f
C582 a_n1236_n9479.n37 vss 0.194658f
C583 a_n1236_n9479.t4 vss 0.428407f
C584 a_n1236_n9479.t0 vss 0.429046f
C585 a_n1236_n9479.t21 vss 0.036678f
C586 a_n1236_n9479.t38 vss 0.036678f
C587 a_n1236_n9479.n38 vss 0.078351f
C588 a_n1236_n9479.t42 vss 0.036678f
C589 a_n1236_n9479.t1 vss 0.036678f
C590 a_n1236_n9479.n39 vss 0.078351f
C591 a_n1236_n9479.n40 vss 0.281102f
C592 a_n1236_n9479.n41 vss 0.512311f
C593 a_n1236_n9479.n42 vss 0.190453f
C594 a_n1236_n9479.t23 vss 0.036678f
C595 a_n1236_n9479.t47 vss 0.036678f
C596 a_n1236_n9479.n43 vss 0.078298f
C597 a_n1236_n9479.t34 vss 0.036678f
C598 a_n1236_n9479.t11 vss 0.036678f
C599 a_n1236_n9479.n44 vss 0.078298f
C600 a_n1236_n9479.n45 vss 0.192954f
C601 a_n1236_n9479.t24 vss 0.428407f
C602 a_n1236_n9479.n46 vss 0.126637f
C603 a_n1236_n9479.n47 vss 0.229843f
C604 a_n1236_n9479.t10 vss 0.428407f
C605 a_n1236_n9479.n48 vss 0.19241f
C606 a_n1236_n9479.n49 vss 0.196776f
C607 a_n1236_n9479.n50 vss 0.133795f
C608 a_n1236_n9479.t25 vss 0.036678f
C609 a_n1236_n9479.t32 vss 0.036678f
C610 a_n1236_n9479.n51 vss 0.078298f
C611 a_n1236_n9479.t43 vss 0.036678f
C612 a_n1236_n9479.t9 vss 0.036678f
C613 a_n1236_n9479.n52 vss 0.078298f
C614 a_n1236_n9479.t27 vss 0.036678f
C615 a_n1236_n9479.t33 vss 0.036678f
C616 a_n1236_n9479.n53 vss 0.078508f
C617 a_n1236_n9479.n54 vss 0.109851f
C618 a_n1236_n9479.n55 vss 0.128037f
C619 a_n1236_n9479.t26 vss 0.428407f
C620 a_n1236_n9479.n56 vss 0.194392f
C621 a_n1236_n9479.n57 vss 0.192707f
C622 a_n1236_n9479.t8 vss 0.428407f
C623 a_n1236_n9479.n58 vss 0.252273f
C624 a_n1236_n9479.n59 vss 0.285147f
C625 a_n1236_n9479.n60 vss 0.138692f
C626 a_n1236_n9479.n61 vss 0.126601f
C627 a_n1236_n9479.n62 vss 0.195682f
C628 a_n1236_n9479.t20 vss 0.428407f
C629 a_n1236_n9479.n63 vss 0.185109f
C630 a_n1236_n9479.n64 vss 0.213178f
C631 a_n1236_n9479.n65 vss 0.126622f
C632 a_n1236_n9479.n66 vss 0.074228f
C633 a_n1236_n9479.t41 vss 0.036678f
C634 a_n1236_n9479.t5 vss 0.036678f
C635 a_n1236_n9479.n67 vss 0.078351f
C636 a_n1236_n9479.n68 vss 0.224594f
C637 a_n1236_n9479.t19 vss 0.036678f
C638 a_n1236_n9479.t44 vss 0.036678f
C639 a_n1236_n9479.n69 vss 0.078351f
C640 a_n1236_n9479.n70 vss 0.191262f
C641 a_n1236_n9479.t18 vss 0.428407f
C642 a_n1236_n9479.n71 vss 0.181786f
C643 a_n1236_n9479.n72 vss 0.116531f
C644 a_n1236_n9479.n73 vss 0.075366f
C645 a_n1236_n9479.n74 vss 0.116443f
C646 a_n1236_n9479.n75 vss 0.160573f
C647 a_n1236_n9479.n76 vss 0.15275f
C648 a_n1236_n9479.n77 vss 0.230436f
C649 a_n1236_n9479.n78 vss 0.126601f
C650 a_n1236_n9479.n79 vss 0.188243f
C651 a_n1236_n9479.t22 vss 0.428407f
C652 a_n1236_n9479.n80 vss 0.192695f
C653 a_n1236_n9479.t12 vss 0.428407f
C654 a_n1236_n9479.n81 vss 0.191841f
C655 a_n1236_n9479.n82 vss 0.126638f
C656 a_n1236_n9479.t35 vss 0.036678f
C657 a_n1236_n9479.t13 vss 0.036678f
C658 a_n1236_n9479.n83 vss 0.078298f
C659 a_n1236_n9479.n84 vss 0.078298f
C660 a_n1236_n9479.t31 vss 0.036678f
C661 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 vss 4.489069f
C662 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 vss 5.32305f
C663 OTA_vref_0.OTA_vref_stage2_0.vref0.t0 vss 0.077096f
C664 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 vss 0.07938f
C665 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 vss 0.07938f
C666 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 vss 0.264281f
C667 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 vss 0.07938f
C668 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 vss 0.07938f
C669 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 vss 0.254416f
C670 OTA_vref_0.OTA_vref_stage2_0.vref0.t32 vss 0.07938f
C671 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 vss 0.07938f
C672 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 vss 0.254416f
C673 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 vss 0.07938f
C674 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 vss 0.07938f
C675 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 vss 0.254416f
C676 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 vss 0.07938f
C677 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 vss 0.07938f
C678 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 vss 0.254416f
C679 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 vss 0.07938f
C680 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 vss 0.07938f
C681 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 vss 0.254416f
C682 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 vss 0.07938f
C683 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 vss 0.07938f
C684 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 vss 0.278065f
C685 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 vss 0.07938f
C686 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 vss 0.07938f
C687 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 vss 0.254416f
C688 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 vss 0.07938f
C689 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 vss 0.07938f
C690 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 vss 0.254416f
C691 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 vss 0.07938f
C692 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 vss 0.07938f
C693 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 vss 0.254416f
C694 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 vss 0.07938f
C695 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 vss 0.07938f
C696 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 vss 0.254416f
C697 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 vss 0.07938f
C698 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 vss 0.07938f
C699 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 vss 0.254416f
C700 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 vss 0.07938f
C701 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 vss 0.07938f
C702 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 vss 0.254416f
C703 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 vss 0.07938f
C704 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 vss 0.07938f
C705 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 vss 0.254416f
C706 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 vss 0.07938f
C707 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 vss 0.07938f
C708 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 vss 0.254284f
C709 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 vss 0.07938f
C710 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 vss 0.07938f
C711 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 vss 0.254416f
C712 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 vss 0.072231f
C713 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 vss 0.110183f
C714 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 vss 0.109159f
C715 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 vss -3.70902f
C716 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 vss 3.98388f
C717 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 vss 0.478981f
C718 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 vss 0.480213f
C719 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 vss 1.17119f
C720 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 vss 0.305431f
C721 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 vss 0.478028f
C722 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 vss 0.234187f
C723 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 vss 0.470573f
C724 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 vss 0.478028f
C725 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 vss 0.470573f
C726 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 vss 0.478028f
C727 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 vss 0.470129f
C728 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 vss 0.478028f
C729 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 vss 0.119324f
C730 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 vss 0.391163f
C731 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 vss 0.207747f
C732 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 vss 0.305316f
C733 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 vss 0.478809f
C734 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 vss 0.222027f
C735 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 vss 0.474153f
C736 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 vss 0.478028f
C737 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 vss 0.474153f
C738 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 vss 0.478028f
C739 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 vss 0.472108f
C740 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 vss 0.478028f
C741 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 vss 0.114607f
C742 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 vss 0.358056f
C743 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 vss 0.1713f
C744 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 vss 0.305164f
C745 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 vss 0.478028f
C746 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 vss 0.234725f
C747 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 vss 0.471116f
C748 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 vss 0.478028f
C749 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 vss 0.471116f
C750 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 vss 0.478028f
C751 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 vss 0.471016f
C752 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 vss 0.478028f
C753 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 vss 0.116651f
C754 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 vss 0.391917f
C755 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 vss 0.175402f
C756 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 vss 0.305187f
C757 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 vss 0.478881f
C758 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 vss 0.232796f
C759 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 vss 0.470031f
C760 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 vss 0.478028f
C761 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 vss 0.470031f
C762 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 vss 0.478028f
C763 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 vss 0.470335f
C764 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 vss 0.478028f
C765 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 vss 0.118954f
C766 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 vss 0.357235f
C767 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 vss 0.171379f
C768 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 vss 0.305728f
C769 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 vss 0.478028f
C770 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 vss 0.231521f
C771 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 vss 0.470851f
C772 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 vss 0.478028f
C773 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 vss 0.470852f
C774 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 vss 0.478028f
C775 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 vss 0.466741f
C776 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 vss 0.478028f
C777 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 vss 0.124091f
C778 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 vss 0.391922f
C779 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 vss 0.175402f
C780 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 vss 0.478028f
C781 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 vss 0.28265f
C782 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 vss 0.46793f
C783 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 vss 0.478028f
C784 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 vss 0.240285f
C785 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 vss 0.478028f
C786 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 vss 0.46793f
C787 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 vss 0.304748f
C788 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 vss 0.478028f
C789 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 vss 0.303889f
C790 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 vss 0.157732f
C791 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 vss 0.205161f
C792 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 vss 0.171854f
C793 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 vss 0.305508f
C794 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 vss 0.478028f
C795 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 vss 0.22844f
C796 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 vss 0.473853f
C797 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 vss 0.478028f
C798 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 vss 0.473853f
C799 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 vss 0.478028f
C800 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 vss 0.473079f
C801 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 vss 0.478028f
C802 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 vss 0.113695f
C803 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 vss 0.395354f
C804 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 vss 0.17643f
C805 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 vss 0.480413f
C806 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 vss 0.478986f
C807 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 vss 1.18519f
C808 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 vss 0.383039f
C809 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 vss 0.473185f
C810 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 vss 0.215214f
C811 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 vss 0.201225f
C812 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 vss 0.215214f
C813 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 vss 0.215214f
C814 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 vss 0.184059f
C815 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 vss 0.04125f
C816 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 vss 0.041255f
C817 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 vss 1.0568f
C818 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 vss 0.444711f
C819 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 vss 0.122425f
C820 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 vss 0.110183f
C821 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 vss 0.10796f
C822 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 vss 0.122425f
C823 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 vss 0.490623f
C824 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 vss 0.201231f
C825 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 vss 0.381488f
C826 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 vss 0.147422f
C827 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 vss 0.329195f
C828 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 vss 0.122425f
C829 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 vss 0.21592f
C830 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 vss 0.21592f
C831 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 vss 0.101613f
C832 a_7434_495.n0 vss 1.46343f
C833 a_7434_495.n1 vss 0.936679f
C834 a_7434_495.n2 vss 1.29294f
C835 a_7434_495.n3 vss 5.4296f
C836 a_7434_495.n4 vss 0.906851f
C837 a_7434_495.n5 vss 0.620305f
C838 a_7434_495.n6 vss 0.742801f
C839 a_7434_495.n7 vss 0.763129f
C840 a_7434_495.n8 vss 1.26286f
C841 a_7434_495.t0 vss 0.150205f
C842 a_7434_495.t12 vss 0.127287f
C843 a_7434_495.t8 vss 1.5052f
C844 a_7434_495.t9 vss 0.080806f
C845 a_7434_495.t10 vss 1.48973f
C846 a_7434_495.t7 vss 0.021976f
C847 a_7434_495.t11 vss 0.021976f
C848 a_7434_495.n9 vss 0.044771f
C849 a_7434_495.t6 vss 1.48363f
C850 a_7434_495.t4 vss 1.49909f
C851 a_7434_495.t5 vss 0.080806f
C852 a_7434_495.t1 vss 0.026371f
C853 a_7434_495.t2 vss 0.026371f
C854 a_7434_495.n10 vss 0.083184f
C855 a_7434_495.t3 vss 0.13999f
C856 2nd_3_OTA_0.vd3.n0 vss 0.456197f
C857 2nd_3_OTA_0.vd3.n1 vss 1.97994f
C858 2nd_3_OTA_0.vd3.n2 vss 1.83635f
C859 2nd_3_OTA_0.vd3.n3 vss 0.036861f
C860 2nd_3_OTA_0.vd3.n4 vss 1.84565f
C861 2nd_3_OTA_0.vd3.n5 vss 2.01845f
C862 2nd_3_OTA_0.vd3.t19 vss 0.292323f
C863 2nd_3_OTA_0.vd3.t18 vss 0.292237f
C864 2nd_3_OTA_0.vd3.t13 vss 0.292237f
C865 2nd_3_OTA_0.vd3.t12 vss 0.291885f
C866 2nd_3_OTA_0.vd3.t2 vss 0.218393f
C867 2nd_3_OTA_0.vd3.t1 vss 0.241422f
C868 2nd_3_OTA_0.vd3.t3 vss 0.047867f
C869 2nd_3_OTA_0.vd3.t0 vss 0.047867f
C870 2nd_3_OTA_0.vd3.n6 vss 0.150893f
C871 2nd_3_OTA_0.vd3.n7 vss 0.638972f
C872 2nd_3_OTA_0.vd3.t11 vss 0.016894f
C873 2nd_3_OTA_0.vd3.t9 vss 0.016894f
C874 2nd_3_OTA_0.vd3.t8 vss 0.665688f
C875 2nd_3_OTA_0.vd3.t16 vss 0.665686f
C876 2nd_3_OTA_0.vd3.n8 vss 0.248119f
C877 2nd_3_OTA_0.vd3.t15 vss 0.665688f
C878 2nd_3_OTA_0.vd3.t4 vss 0.665686f
C879 2nd_3_OTA_0.vd3.n9 vss 0.248119f
C880 2nd_3_OTA_0.vd3.t5 vss 0.004787f
C881 2nd_3_OTA_0.vd3.t7 vss 0.004787f
C882 2nd_3_OTA_0.vd3.n10 vss 0.010125f
C883 2nd_3_OTA_0.vd3.t17 vss 0.665688f
C884 2nd_3_OTA_0.vd3.t6 vss 0.665686f
C885 2nd_3_OTA_0.vd3.n11 vss 0.248119f
C886 2nd_3_OTA_0.vd3.t10 vss 0.665688f
C887 2nd_3_OTA_0.vd3.t14 vss 0.665686f
C888 2nd_3_OTA_0.vd3.n12 vss 0.248119f
C889 2nd_3_OTA_0.vd3.n13 vss 1.78256f
.ends

