magic
tech sky130A
magscale 1 2
timestamp 1738105933
<< nwell >>
rect 11101 1517 19111 2992
<< pwell >>
rect 12365 -2528 17892 1027
rect 12449 -2562 12472 -2528
rect 12566 -2562 17799 -2560
<< psubdiff >>
rect 12418 940 12478 974
rect 17779 940 17839 974
rect 12418 914 12452 940
rect 17805 914 17839 940
rect 12418 -2454 12452 -2428
rect 17805 -2454 17839 -2428
rect 12418 -2488 12478 -2454
rect 17779 -2488 17839 -2454
<< nsubdiff >>
rect 11187 2901 11247 2935
rect 18935 2901 18995 2935
rect 11187 2875 11221 2901
rect 11187 1593 11221 1619
rect 18961 2875 18995 2901
rect 18961 1593 18995 1619
rect 11187 1559 11247 1593
rect 18935 1559 18995 1593
<< psubdiffcont >>
rect 12478 940 17779 974
rect 12418 -2428 12452 914
rect 17805 -2428 17839 914
rect 12478 -2488 17779 -2454
<< nsubdiffcont >>
rect 11247 2901 18935 2935
rect 11187 1619 11221 2875
rect 18961 1619 18995 2875
rect 11247 1559 18935 1593
<< poly >>
rect 14674 -2388 14821 -2336
<< locali >>
rect 10995 3080 19171 3116
rect 10995 2991 11179 3080
rect 18977 2991 19171 3080
rect 10995 2935 19171 2991
rect 10995 2901 11247 2935
rect 18935 2901 19171 2935
rect 10995 2875 19171 2901
rect 10995 1619 11187 2875
rect 11221 2778 18961 2875
rect 11221 1619 11249 2778
rect 10995 1609 11249 1619
rect 18995 2778 19171 2875
rect 18995 1619 19170 2778
rect 18961 1609 19170 1619
rect 10995 1593 19170 1609
rect 10995 1559 11247 1593
rect 18935 1559 19170 1593
rect 10995 1476 19170 1559
rect 10996 974 18145 1041
rect 10996 940 12478 974
rect 17779 940 18145 974
rect 10996 914 18145 940
rect 10996 -640 12418 914
rect 10995 -677 12418 -640
rect 10995 -1923 11206 -677
rect 11311 -1923 11919 -1841
rect 12047 -1923 12418 -677
rect 10995 -2153 12418 -1923
rect 10993 -2357 12418 -2153
rect 10993 -2451 11101 -2357
rect 11654 -2428 12418 -2357
rect 12452 901 17805 914
rect 12452 -2428 12472 901
rect 11654 -2433 12472 -2428
rect 17795 -2428 17805 901
rect 17839 -2428 18145 914
rect 17795 -2433 18145 -2428
rect 11654 -2451 18145 -2433
rect 10993 -2454 18145 -2451
rect 10993 -2488 12478 -2454
rect 17779 -2488 18145 -2454
rect 10993 -2592 18145 -2488
rect 10993 -2681 11103 -2592
rect 18037 -2681 18145 -2592
rect 10993 -2743 18145 -2681
<< viali >>
rect 11179 2991 18977 3080
rect 11101 -2451 11654 -2357
rect 11103 -2681 18037 -2592
<< metal1 >>
rect 11167 3080 18989 3086
rect 11167 2991 11179 3080
rect 18977 2991 18989 3080
rect 11167 2985 18989 2991
rect 11297 2281 11497 2729
rect 11297 1250 11383 2281
rect 11411 2111 11497 2154
rect 11487 1806 11497 2111
rect 11411 1793 11497 1806
rect 11674 1751 14913 2696
rect 15074 2683 15190 2729
rect 15082 2294 15092 2630
rect 15146 2294 15156 2630
rect 15082 1806 15092 2142
rect 15146 1806 15156 2142
rect 15050 1707 15166 1753
rect 15336 1751 18575 2696
rect 18740 2283 18942 2643
rect 18742 2101 18828 2154
rect 18742 1806 18752 2101
rect 18742 1707 18828 1806
rect 18856 1435 18942 2283
rect 11411 1428 19170 1435
rect 11720 1420 19170 1428
rect 11720 1353 12219 1420
rect 12568 1417 19170 1420
rect 12568 1353 17283 1417
rect 11720 1350 17283 1353
rect 17632 1350 19170 1417
rect 11720 1344 19170 1350
rect 11411 1335 19170 1344
rect 11297 1234 18838 1250
rect 11297 1230 17703 1234
rect 11297 1163 12646 1230
rect 12995 1167 17703 1230
rect 18052 1167 18417 1234
rect 12995 1164 18417 1167
rect 18807 1164 18838 1234
rect 12995 1163 18838 1164
rect 11297 1150 18838 1163
rect 12600 190 12610 758
rect 12696 190 12706 758
rect 12600 -376 12706 190
rect 13352 -456 14437 813
rect 15094 -386 15104 -67
rect 15156 -386 15166 -67
rect 15856 -456 16943 808
rect 17552 190 17562 758
rect 17648 190 17658 758
rect 17552 -363 17658 190
rect 12710 -513 12720 -456
rect 12930 -513 15094 -456
rect 15164 -513 17332 -456
rect 17542 -513 17552 -456
rect 12720 -574 15173 -570
rect 12720 -631 12743 -574
rect 12930 -631 15173 -574
rect 12720 -634 15173 -631
rect 15374 -634 15383 -570
rect 12720 -649 15383 -634
rect 11317 -793 11327 -738
rect 11903 -793 11913 -738
rect 11947 -986 12006 -805
rect 14873 -887 17542 -867
rect 14873 -889 17332 -887
rect 15083 -944 17332 -889
rect 15083 -946 17542 -944
rect 14873 -956 17542 -946
rect 11935 -1004 11945 -986
rect 11279 -1601 11945 -1004
rect 11935 -1785 11945 -1601
rect 11997 -1785 12007 -986
rect 12705 -1078 14873 -1021
rect 15083 -1078 15093 -1021
rect 11947 -1797 12006 -1785
rect 12494 -2189 12543 -1117
rect 12695 -2189 12705 -1117
rect 12494 -2258 12705 -2189
rect 13347 -2336 14434 -1078
rect 15163 -1079 15173 -1022
rect 15383 -1079 17551 -1022
rect 15093 -1467 15103 -1148
rect 15155 -1467 15165 -1148
rect 11089 -2357 11666 -2351
rect 11089 -2451 11101 -2357
rect 11654 -2451 11666 -2357
rect 12703 -2388 12715 -2336
rect 13195 -2388 15095 -2336
rect 15163 -2387 15173 -2335
rect 15653 -2387 15663 -2335
rect 15847 -2337 16934 -1079
rect 17550 -2189 17560 -1117
rect 17712 -2189 17722 -1117
rect 11089 -2457 11666 -2451
rect 11091 -2592 18049 -2586
rect 11091 -2681 11103 -2592
rect 18037 -2681 18049 -2592
rect 11091 -2687 18049 -2681
<< via1 >>
rect 11179 2991 18977 3080
rect 11411 1806 11487 2111
rect 15092 2294 15146 2630
rect 15092 1806 15146 2142
rect 18752 1806 18828 2101
rect 11411 1344 11720 1428
rect 12219 1353 12568 1420
rect 17283 1350 17632 1417
rect 12646 1163 12995 1230
rect 17703 1167 18052 1234
rect 18417 1164 18807 1234
rect 12610 190 12696 758
rect 15104 -386 15156 -67
rect 17562 190 17648 758
rect 12720 -513 12930 -456
rect 17332 -513 17542 -456
rect 12743 -631 12930 -574
rect 15173 -634 15374 -570
rect 11327 -793 11903 -738
rect 14873 -946 15083 -889
rect 17332 -944 17542 -887
rect 11945 -1785 11997 -986
rect 14873 -1078 15083 -1021
rect 12543 -2189 12695 -1117
rect 15173 -1079 15383 -1022
rect 15103 -1467 15155 -1148
rect 11101 -2451 11654 -2357
rect 12715 -2388 13195 -2336
rect 15173 -2387 15653 -2335
rect 17560 -2189 17712 -1117
rect 11103 -2681 18037 -2592
<< metal2 >>
rect 10995 3080 19171 3381
rect 10995 2991 11179 3080
rect 18977 2991 19171 3080
rect 10995 2981 19171 2991
rect 15092 2630 15146 2981
rect 11401 2111 11487 2154
rect 11401 1806 11411 2111
rect 11401 1438 11487 1806
rect 15092 2142 15146 2294
rect 15092 1796 15146 1806
rect 18752 2101 18838 2154
rect 18828 1806 18838 2101
rect 11401 1428 11720 1438
rect 11401 1344 11411 1428
rect 11401 1334 11720 1344
rect 12219 1420 12580 1435
rect 12568 1353 12580 1420
rect 12219 1335 12580 1353
rect 17283 1417 17648 1435
rect 17632 1350 17648 1417
rect 17283 1335 17648 1350
rect 11327 -728 11903 -718
rect 11327 -803 11903 -793
rect 11945 -977 11997 -976
rect 11942 -986 12000 -977
rect 11942 -987 11945 -986
rect 11997 -987 12000 -986
rect 11942 -1795 12000 -1785
rect 12494 -1107 12580 1335
rect 12610 1230 12996 1250
rect 12610 1163 12646 1230
rect 12995 1163 12996 1230
rect 12610 1150 12996 1163
rect 12610 758 12696 1150
rect 12610 180 12696 190
rect 17562 758 17648 1335
rect 18752 1250 18838 1806
rect 17562 180 17648 190
rect 17678 1234 18052 1250
rect 17678 1167 17703 1234
rect 17678 1150 18052 1167
rect 18417 1234 18838 1250
rect 18807 1164 18838 1234
rect 18417 1150 18838 1164
rect 15100 -54 15156 -44
rect 15100 -406 15156 -396
rect 12720 -456 12930 -446
rect 12720 -574 12930 -513
rect 17332 -456 17542 -446
rect 12720 -631 12743 -574
rect 12720 -641 12930 -631
rect 15173 -570 15383 -558
rect 15374 -634 15383 -570
rect 14873 -889 15083 -879
rect 14873 -1021 15083 -946
rect 14873 -1088 15083 -1078
rect 15173 -1022 15383 -634
rect 17332 -887 17542 -513
rect 17332 -954 17542 -944
rect 15173 -1089 15383 -1079
rect 17678 -1107 17764 1150
rect 12494 -1117 12695 -1107
rect 12494 -2189 12543 -1117
rect 17560 -1117 17764 -1107
rect 15099 -1138 15157 -1128
rect 15099 -1487 15157 -1477
rect 12695 -2189 12697 -1681
rect 12494 -2258 12697 -2189
rect 17712 -2189 17764 -1117
rect 17560 -2199 17764 -2189
rect 10993 -2357 11775 -2291
rect 10993 -2451 11101 -2357
rect 11654 -2451 11775 -2357
rect 12715 -2333 13195 -2323
rect 12715 -2401 13195 -2391
rect 15173 -2331 15653 -2321
rect 15173 -2399 15653 -2389
rect 10993 -2582 11775 -2451
rect 10993 -2592 18037 -2582
rect 10993 -2681 11103 -2592
rect 10993 -2691 18037 -2681
<< via2 >>
rect 11327 -738 11903 -728
rect 11327 -793 11903 -738
rect 11942 -1785 11945 -987
rect 11945 -1785 11997 -987
rect 11997 -1785 12000 -987
rect 15100 -67 15156 -54
rect 15100 -386 15104 -67
rect 15104 -386 15156 -67
rect 15100 -396 15156 -386
rect 15099 -1148 15157 -1138
rect 15099 -1467 15103 -1148
rect 15103 -1467 15155 -1148
rect 15155 -1467 15157 -1148
rect 15099 -1477 15157 -1467
rect 12715 -2336 13195 -2333
rect 12715 -2388 13195 -2336
rect 12715 -2391 13195 -2388
rect 15173 -2335 15653 -2331
rect 15173 -2387 15653 -2335
rect 15173 -2389 15653 -2387
<< metal3 >>
rect 15089 -54 15167 -49
rect 15089 -396 15100 -54
rect 15156 -396 15167 -54
rect 15089 -723 15167 -396
rect 11317 -728 15167 -723
rect 11317 -793 11327 -728
rect 11903 -793 15167 -728
rect 11317 -798 15167 -793
rect 11932 -987 12112 -982
rect 11932 -1785 11942 -987
rect 12000 -1785 12112 -987
rect 15089 -1138 15167 -798
rect 15089 -1477 15099 -1138
rect 15157 -1477 15167 -1138
rect 15089 -1482 15167 -1477
rect 11932 -2832 12112 -1785
rect 12705 -2333 13205 -2328
rect 12705 -2391 12715 -2333
rect 13195 -2391 13205 -2333
rect 12705 -2396 13205 -2391
rect 15163 -2331 15663 -2326
rect 15163 -2389 15173 -2331
rect 15653 -2389 15663 -2331
rect 15163 -2394 15663 -2389
rect 12705 -2832 12885 -2396
rect 15163 -2828 15343 -2394
use sky130_fd_pr__nfet_01v8_lvt_59CFV9  sky130_fd_pr__nfet_01v8_lvt_59CFV9_0
timestamp 1737073392
transform 1 0 16358 0 1 170
box -1258 -688 1258 688
use sky130_fd_pr__pfet_01v8_lvt_58FN7G  sky130_fd_pr__pfet_01v8_lvt_58FN7G_0
timestamp 1737085049
transform 1 0 16948 0 1 2462
box -1894 -280 1894 280
use sky130_fd_pr__nfet_01v8_lvt_59CFV9  XM1
timestamp 1737073392
transform 1 0 13900 0 1 170
box -1258 -688 1258 688
use sky130_fd_pr__nfet_01v8_lvt_59CFV9  XM2
timestamp 1737073392
transform 1 0 13899 0 1 -1705
box -1258 -688 1258 688
use sky130_fd_pr__nfet_01v8_Q93DRV  XM3
timestamp 1737072185
transform 0 -1 11615 1 0 -1301
box -696 -510 696 510
use sky130_fd_pr__pfet_01v8_lvt_58FN7G  XM4
timestamp 1737085049
transform 1 0 13290 0 -1 1974
box -1894 -280 1894 280
use sky130_fd_pr__pfet_01v8_lvt_58FN7G  XM5
timestamp 1737085049
transform 1 0 13290 0 -1 2462
box -1894 -280 1894 280
use sky130_fd_pr__pfet_01v8_lvt_58FN7G  XM6
timestamp 1737085049
transform 1 0 16948 0 1 1974
box -1894 -280 1894 280
use sky130_fd_pr__nfet_01v8_lvt_59CFV9  XM8
timestamp 1737073392
transform 1 0 16357 0 1 -1705
box -1258 -688 1258 688
<< labels >>
rlabel metal1 19169 1388 19169 1388 3 vout
port 1 e
rlabel metal3 15247 -2825 15247 -2825 5 vin_p
port 2 s
rlabel metal3 12781 -2829 12781 -2829 5 vin_n
port 3 s
rlabel metal3 12014 -2831 12014 -2831 5 vb
port 4 s
rlabel metal2 10996 3203 10996 3203 7 vcc
port 5 w
rlabel metal2 10994 -2533 10994 -2533 7 vss
port 6 w
<< end >>
