* NGSPICE file created from BGR_BJT_stage1.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2 a_100_n400# a_n158_n400# a_n100_n488# VSUBS
X0 a_100_n400# a_n100_n488# a_n158_n400# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_QCPJZY a_n100_n197# a_100_n100# w_n194_n200# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n194_n200# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_KLHH7J a_n200_n147# a_n258_n50# a_200_n50# w_n294_n150#
X0 a_200_n50# a_n200_n147# a_n258_n50# w_n294_n150# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
.ends

.subckt BGR_BJT_stage1 vcc vss vref0 vr
XXM12 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM23 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM34 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM45 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM25 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM24 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM36 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM35 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM47 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM46 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM14 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM26 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM37 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM48 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM15 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM27 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM38 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM49 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM16 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM28 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM39 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM17 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM18 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM29 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM19 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM1 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM2 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM3 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM4 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM5 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM6 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM7 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM9 vr vcc vcc sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter sky130_fd_pr__pfet_01v8_lvt_QCPJZY
XXM8 vr vr vcc vcc sky130_fd_pr__pfet_01v8_lvt_KLHH7J
Xsky130_fd_pr__nfet_01v8_lvt_UZ3GQ2_0 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM50 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__pfet_01v8_lvt_KLHH7J_0 vr vcc vr vcc sky130_fd_pr__pfet_01v8_lvt_KLHH7J
XXM40 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__pfet_01v8_lvt_QCPJZY_0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
+ vcc vcc sky130_fd_pr__pfet_01v8_lvt_QCPJZY
XXM41 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM30 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
+ vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXM42 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM20 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM31 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM10 vr vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM21 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM32 m1_9688_899# vref0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM43 m1_9688_899# vss m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM11 vref0 vr sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM22 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM33 vref0 m1_9688_899# sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
XXM44 vss m1_9688_899# m1_9688_899# vss sky130_fd_pr__nfet_01v8_lvt_UZ3GQ2
.ends

