magic
tech sky130A
magscale 1 2
timestamp 1741310630
<< nwell >>
rect -820 484 4074 2918
<< pwell >>
rect 556 3053 2692 5338
<< psubdiff >>
rect 572 5279 632 5313
rect 2614 5279 2674 5313
rect 572 5253 606 5279
rect 572 3109 606 3135
rect 2640 5253 2674 5279
rect 3748 4766 3808 4800
rect 4407 4766 4467 4800
rect 3748 4740 3782 4766
rect 3748 4274 3782 4300
rect 4433 4740 4467 4766
rect 4433 4274 4467 4300
rect 3748 4240 3808 4274
rect 4407 4240 4467 4274
rect 2640 3109 2674 3135
rect 572 3075 632 3109
rect 2614 3075 2674 3109
<< nsubdiff >>
rect -768 2827 -708 2861
rect 3978 2827 4038 2861
rect -768 2801 -734 2827
rect -768 562 -734 588
rect 4004 2801 4038 2827
rect 4004 562 4038 588
rect -768 528 -708 562
rect 3978 528 4038 562
<< psubdiffcont >>
rect 632 5279 2614 5313
rect 572 3135 606 5253
rect 2640 3135 2674 5253
rect 3808 4766 4407 4800
rect 3748 4300 3782 4740
rect 4433 4300 4467 4740
rect 3808 4240 4407 4274
rect 632 3075 2614 3109
<< nsubdiffcont >>
rect -708 2827 3978 2861
rect -768 588 -734 2801
rect 4004 588 4038 2801
rect -708 528 3978 562
<< locali >>
rect 494 6770 2647 6821
rect 494 6761 2392 6770
rect 494 5571 503 6761
rect 730 6759 2392 6761
rect 491 5334 503 5571
rect 841 6441 2392 6520
rect 841 5571 977 6441
rect 2335 5571 2392 6441
rect 841 5504 2392 5571
rect 2603 5571 2647 6770
rect 2720 5571 4559 5572
rect 2603 5508 4559 5571
rect 2603 5504 3210 5508
rect 491 5233 548 5334
rect 622 5313 2630 5334
rect 622 5279 632 5313
rect 2614 5279 2630 5313
rect 537 4703 548 5233
rect 622 5233 2630 5279
rect 622 4703 630 5233
rect 537 3667 572 4703
rect 606 3667 630 4703
rect 537 3151 557 3667
rect 530 3026 557 3151
rect 615 3151 630 3667
rect 2617 3151 2630 5233
rect 615 3129 2630 3151
rect 2706 5232 3048 5334
rect 2706 3123 2739 5232
rect 3025 4886 3048 5232
rect 3168 5296 3210 5504
rect 4488 5296 4559 5508
rect 3168 5158 4559 5296
rect 4426 4886 4559 5158
rect 3025 4800 4559 4886
rect 3025 4766 3808 4800
rect 4407 4766 4559 4800
rect 3025 4749 4559 4766
rect 3025 4740 3800 4749
rect 3025 4300 3748 4740
rect 3782 4300 3800 4740
rect 3025 4298 3800 4300
rect 4413 4740 4559 4749
rect 4413 4300 4433 4740
rect 4467 4300 4559 4740
rect 4413 4298 4559 4300
rect 3025 4274 4559 4298
rect 3025 4240 3808 4274
rect 4407 4240 4559 4274
rect 3025 4220 4559 4240
rect 3623 4052 3761 4135
rect 2706 3026 2731 3123
rect 530 3001 2731 3026
rect 3623 2920 3644 4052
rect -808 2914 3644 2920
rect -822 2893 3644 2914
rect 3748 3279 3761 4052
rect 4424 3279 4507 4121
rect -822 2886 -766 2893
rect -822 706 -801 2886
rect 3748 2861 4507 3279
rect 3978 2838 4507 2861
rect 3978 2827 4120 2838
rect 3748 2801 4120 2827
rect -1013 594 -801 706
rect -1013 229 -863 594
rect 3748 2796 4004 2801
rect -684 2762 4004 2796
rect -684 706 -642 2762
rect 3962 1407 4004 2762
rect 4038 1407 4120 2801
rect 3962 706 3983 1407
rect -684 594 3983 706
rect 3941 593 3983 594
rect 4080 593 4120 1407
rect 4099 560 4120 593
rect -1013 228 3840 229
rect 4099 228 4117 560
rect -1013 -144 4117 228
<< viali >>
rect 503 6759 730 6761
rect 2392 6759 2603 6770
rect 503 6520 2603 6759
rect 503 5504 841 6520
rect 2392 5504 2603 6520
rect 503 5334 3168 5504
rect 548 5253 622 5334
rect 548 4703 572 5253
rect 572 4703 606 5253
rect 606 4703 622 5253
rect 2630 5253 2706 5334
rect 557 3135 572 3667
rect 572 3135 606 3667
rect 606 3135 615 3667
rect 557 3129 615 3135
rect 2630 3135 2640 5253
rect 2640 3135 2674 5253
rect 2674 3135 2706 5253
rect 2630 3129 2706 3135
rect 557 3109 2706 3129
rect 3048 5158 3168 5334
rect 3048 4886 4426 5158
rect 557 3075 632 3109
rect 632 3075 2614 3109
rect 2614 3075 2706 3109
rect 557 3026 2706 3075
rect 3644 2893 3748 4052
rect -766 2886 3748 2893
rect -801 2861 3748 2886
rect -801 2827 -708 2861
rect -708 2827 3748 2861
rect -801 2801 3748 2827
rect -801 594 -768 2801
rect -863 588 -768 594
rect -768 588 -734 2801
rect -734 2796 3748 2801
rect -734 594 -684 2796
rect -734 593 3941 594
rect 3983 593 4004 1407
rect -734 588 4004 593
rect 4004 588 4038 1407
rect 4038 593 4080 1407
rect 4038 588 4099 593
rect -863 562 4099 588
rect -863 528 -708 562
rect -708 528 3978 562
rect 3978 528 4099 562
rect -863 229 4099 528
rect 3840 228 4099 229
<< metal1 >>
rect 497 6765 736 6773
rect 2386 6770 2609 6782
rect 2382 6765 2392 6770
rect 497 6761 2392 6765
rect 493 5334 503 6761
rect 730 6759 2392 6761
rect 841 6514 2392 6520
rect 841 5511 851 6514
rect 1760 6336 1770 6401
rect 2179 6336 2189 6401
rect 1053 6120 2228 6281
rect 1013 5976 1059 6047
rect 1093 5979 1103 6043
rect 1603 5979 1613 6043
rect 2223 5976 2269 6046
rect 1053 5853 2228 5926
rect 998 5713 1008 5853
rect 1064 5765 2228 5853
rect 1064 5713 1074 5765
rect 1760 5620 1770 5685
rect 2179 5620 2189 5685
rect 1846 5510 1856 5511
rect 2382 5510 2392 6514
rect 1846 5504 2392 5510
rect 2603 5510 2613 6770
rect 2973 5510 3174 5516
rect 2603 5504 3174 5510
rect 497 5322 548 5334
rect 538 4703 548 5322
rect 622 5328 2630 5334
rect 622 5322 736 5328
rect 622 4703 632 5322
rect 542 4691 628 4703
rect 641 4521 651 4658
rect 745 4521 755 4658
rect 810 4469 1031 5132
rect 1121 4926 1131 5086
rect 1183 4926 1193 5086
rect 1273 4469 1494 5135
rect 1558 4732 1568 4869
rect 1662 4732 1672 4869
rect 1718 4469 1939 5135
rect 2037 4926 2047 5086
rect 2099 4926 2109 5086
rect 2188 4469 2409 5134
rect 2473 4521 2483 4658
rect 2577 4521 2587 4658
rect 734 4417 744 4469
rect 944 4463 1031 4469
rect 944 4417 954 4463
rect 1192 4417 1202 4469
rect 1402 4466 1494 4469
rect 1402 4417 1412 4466
rect 1650 4417 1660 4469
rect 1860 4466 1939 4469
rect 1860 4417 1870 4466
rect 2108 4417 2118 4469
rect 2318 4465 2409 4469
rect 2318 4417 2328 4465
rect -67 4230 744 4330
rect 844 4230 1470 4330
rect 1570 4230 1928 4330
rect 2028 4230 2118 4330
rect 2218 4230 2531 4330
rect -67 4044 1012 4144
rect 1112 4044 1202 4144
rect 1302 4044 1660 4144
rect 1760 4044 2386 4144
rect 2486 4044 2531 4144
rect 902 3926 912 3972
rect 808 3920 912 3926
rect 1112 3920 1122 3972
rect 1360 3926 1370 3972
rect 1267 3920 1370 3926
rect 1570 3920 1580 3972
rect 1818 3926 1828 3972
rect 1730 3920 1828 3926
rect 2028 3920 2038 3972
rect 2276 3925 2286 3972
rect 2184 3920 2286 3925
rect 2486 3920 2496 3972
rect 640 3732 650 3869
rect 744 3732 754 3869
rect 551 3667 621 3679
rect 547 3026 557 3667
rect 615 3135 625 3667
rect 808 3257 1029 3920
rect 1121 3303 1131 3463
rect 1183 3303 1193 3463
rect 1267 3257 1488 3920
rect 1559 3474 1569 3611
rect 1663 3474 1673 3611
rect 1730 3257 1951 3920
rect 2037 3303 2047 3463
rect 2099 3303 2109 3463
rect 2184 3256 2405 3920
rect 2475 3732 2485 3869
rect 2579 3732 2589 3869
rect 2624 3135 2630 5328
rect 615 3129 2630 3135
rect 2706 5328 3048 5334
rect 2706 3026 2712 5328
rect 2973 5322 3048 5328
rect 3042 5164 3048 5322
rect 3036 4886 3048 5164
rect 3168 5164 3174 5504
rect 3334 5378 3344 5430
rect 3546 5378 3556 5430
rect 4168 5379 4178 5431
rect 4380 5379 4390 5431
rect 3168 5158 4438 5164
rect 4426 4886 4438 5158
rect 3036 4880 4438 4886
rect 3942 4646 4311 4692
rect 3851 4531 3861 4602
rect 3913 4531 3923 4602
rect 4207 4531 4217 4602
rect 4269 4531 4279 4602
rect 4295 4426 4305 4497
rect 4357 4426 4367 4497
rect 3958 4382 3992 4419
rect 3939 4303 3949 4382
rect 4001 4336 4269 4382
rect 4001 4303 4011 4336
rect 3638 4052 3754 4064
rect 551 3020 2712 3026
rect 551 3014 621 3020
rect 2624 3014 2712 3020
rect 3634 2899 3644 4052
rect -778 2898 3644 2899
rect -807 2893 3644 2898
rect 3748 2899 3758 4052
rect 3878 3969 3943 4027
rect 4236 3970 4298 4041
rect 3939 3717 3949 3917
rect 4001 3717 4011 3917
rect 4295 3717 4305 3917
rect 4357 3717 4367 3917
rect 3811 3421 3821 3621
rect 3873 3421 3883 3621
rect 4167 3421 4177 3621
rect 4229 3421 4239 3621
rect -807 2886 -766 2893
rect -811 600 -801 2886
rect 3748 2796 3760 2899
rect -875 594 -801 600
rect -684 2790 3760 2796
rect -684 600 -674 2790
rect -509 2547 -452 2593
rect -509 2504 -463 2547
rect -528 2018 -518 2218
rect -454 2018 -444 2218
rect -509 1969 -463 2007
rect -509 1968 -431 1969
rect -271 1968 382 2553
rect 536 2194 546 2494
rect 598 2194 608 2494
rect 761 1968 1414 2552
rect 1594 2547 1665 2593
rect 1607 2506 1653 2547
rect 1588 2294 1598 2494
rect 1662 2294 1672 2494
rect -509 1916 -441 1968
rect 199 1964 382 1968
rect 199 1916 209 1964
rect 607 1916 617 1968
rect 1257 1963 1414 1968
rect 1607 1968 1653 2008
rect 1872 1968 2525 2552
rect 2652 2194 2662 2494
rect 2714 2194 2724 2494
rect 2910 1968 3563 2552
rect 3709 2547 3769 2593
rect 3723 2505 3769 2547
rect 3704 2018 3714 2218
rect 3778 2018 3788 2218
rect 1607 1965 1675 1968
rect 1257 1916 1267 1963
rect 1596 1919 1675 1965
rect 1665 1916 1675 1919
rect 2315 1963 2525 1968
rect 2315 1916 2325 1963
rect 2723 1916 2733 1968
rect 3373 1963 3563 1968
rect 3723 1965 3769 2008
rect 3373 1916 3383 1963
rect 3694 1919 3769 1965
rect -509 1915 -463 1916
rect 3861 1812 3961 3368
rect -457 1712 -441 1812
rect -341 1712 1485 1812
rect 1585 1712 2543 1812
rect 2643 1712 2733 1812
rect 2833 1712 3961 1812
rect 4216 1630 4316 3368
rect -460 1530 427 1630
rect 527 1530 617 1630
rect 717 1530 1675 1630
rect 1775 1530 3601 1630
rect 3701 1530 4316 1630
rect -509 1385 -452 1431
rect -123 1388 -113 1434
rect -509 1343 -463 1385
rect -308 1382 -113 1388
rect 527 1382 537 1434
rect 935 1390 945 1434
rect 778 1382 945 1390
rect 1585 1382 1668 1434
rect 1993 1390 2003 1433
rect -528 1132 -518 1332
rect -454 1132 -444 1332
rect -509 803 -463 851
rect -509 757 -444 803
rect -308 799 345 1382
rect 536 856 546 1156
rect 598 856 608 1156
rect 778 801 1431 1382
rect 1607 1344 1653 1382
rect 1848 1381 2003 1390
rect 2643 1381 2653 1433
rect 3051 1391 3061 1434
rect 2881 1382 3061 1391
rect 3701 1382 3711 1434
rect 3977 1407 4086 1419
rect 1588 856 1598 1056
rect 1662 856 1672 1056
rect 1607 803 1653 846
rect 1596 757 1665 803
rect 1848 801 2501 1381
rect 2652 856 2662 1156
rect 2714 856 2724 1156
rect 2881 802 3534 1382
rect 3704 1132 3714 1332
rect 3778 1132 3788 1332
rect 3723 803 3769 847
rect 3701 757 3769 803
rect 3973 605 3983 1407
rect 3834 600 3983 605
rect -684 594 3983 600
rect -875 229 -863 594
rect 3941 593 3983 594
rect 4080 605 4090 1407
rect 4080 593 4105 605
rect -875 228 3840 229
rect 4099 228 4109 593
rect -875 223 4105 228
rect 3834 216 4105 223
<< via1 >>
rect 503 6759 730 6761
rect 2392 6759 2603 6770
rect 503 6520 2603 6759
rect 503 5504 841 6520
rect 1770 6336 2179 6401
rect 1103 5979 1603 6043
rect 1008 5713 1064 5853
rect 1770 5620 2179 5685
rect 841 5504 1846 5511
rect 503 5341 1846 5504
rect 2392 5469 2603 6520
rect 503 5334 730 5341
rect 548 4703 622 5334
rect 651 4521 745 4658
rect 1131 4926 1183 5086
rect 1568 4732 1662 4869
rect 2047 4926 2099 5086
rect 2483 4521 2577 4658
rect 744 4417 944 4469
rect 1202 4417 1402 4469
rect 1660 4417 1860 4469
rect 2118 4417 2318 4469
rect 744 4230 844 4330
rect 1470 4230 1570 4330
rect 1928 4230 2028 4330
rect 2118 4230 2218 4330
rect 1012 4044 1112 4144
rect 1202 4044 1302 4144
rect 1660 4044 1760 4144
rect 2386 4044 2486 4144
rect 912 3920 1112 3972
rect 1370 3920 1570 3972
rect 1828 3920 2028 3972
rect 2286 3920 2486 3972
rect 650 3732 744 3869
rect 557 3129 615 3667
rect 1131 3303 1183 3463
rect 1569 3474 1663 3611
rect 2047 3303 2099 3463
rect 2485 3732 2579 3869
rect 557 3026 2685 3129
rect 3344 5378 3546 5430
rect 4178 5379 4380 5431
rect 3048 4886 4426 5158
rect 3861 4531 3913 4602
rect 4217 4531 4269 4602
rect 4305 4426 4357 4497
rect 3949 4303 4001 4382
rect 3644 2893 3748 4052
rect 3949 3717 4001 3917
rect 4305 3717 4357 3917
rect 3821 3421 3873 3621
rect 4177 3421 4229 3621
rect -766 2886 3748 2893
rect -801 2796 3748 2886
rect -801 594 -684 2796
rect -518 2018 -454 2218
rect 546 2194 598 2494
rect 1598 2294 1662 2494
rect -441 1916 199 1968
rect 617 1916 1257 1968
rect 2662 2194 2714 2494
rect 3714 2018 3778 2218
rect 1675 1916 2315 1968
rect 2733 1916 3373 1968
rect -441 1712 -341 1812
rect 1485 1712 1585 1812
rect 2543 1712 2643 1812
rect 2733 1712 2833 1812
rect 427 1530 527 1630
rect 617 1530 717 1630
rect 1675 1530 1775 1630
rect 3601 1530 3701 1630
rect -113 1382 527 1434
rect 945 1382 1585 1434
rect -518 1132 -454 1332
rect 546 856 598 1156
rect 2003 1381 2643 1433
rect 3061 1382 3701 1434
rect 1598 856 1662 1056
rect 2662 856 2714 1156
rect 3714 1132 3778 1332
rect -863 593 3941 594
rect 3983 593 4080 1407
rect -863 229 4099 593
rect 3840 228 4099 229
<< metal2 >>
rect 461 6771 621 6772
rect 461 6769 730 6771
rect 2392 6770 2603 6780
rect 461 6761 2392 6769
rect 461 6487 503 6761
rect 730 6759 2392 6761
rect 841 6510 2392 6520
rect 1770 6401 2179 6411
rect 1770 6326 2179 6336
rect 841 6043 1603 6053
rect 841 5979 1103 6043
rect 841 5969 1603 5979
rect 1008 5853 1064 5863
rect 1008 5703 1064 5713
rect 2056 5695 2178 6326
rect 1770 5685 2179 5695
rect 1770 5610 2179 5620
rect 841 5511 1846 5521
rect 730 5334 1846 5341
rect 503 5324 548 5334
rect 622 5331 1846 5334
rect 622 5324 730 5331
rect 2056 5096 2178 5610
rect 2392 5459 2603 5469
rect 3138 5430 3279 5440
rect 3344 5430 3546 5440
rect 3279 5378 3344 5430
rect 3279 5368 3546 5378
rect 4178 5431 4660 5441
rect 4380 5379 4660 5431
rect 4178 5369 4660 5379
rect 3138 5358 3279 5368
rect 1131 5093 1183 5096
rect 2047 5093 2178 5096
rect 3048 5158 4426 5168
rect 1131 5086 2979 5093
rect 1183 4993 2047 5086
rect 1131 4916 1183 4926
rect 2099 4993 2979 5086
rect 2047 4916 2099 4926
rect 1568 4869 1662 4879
rect 1568 4722 1662 4732
rect 548 4693 622 4703
rect 651 4658 745 4668
rect 651 4511 745 4521
rect 2483 4658 2577 4668
rect 2483 4511 2577 4521
rect 744 4469 944 4479
rect 744 4407 944 4417
rect 1202 4469 1402 4479
rect 1202 4407 1402 4417
rect 1660 4469 1860 4479
rect 1660 4407 1860 4417
rect 2118 4469 2318 4479
rect 2118 4407 2318 4417
rect 744 4330 844 4407
rect 744 4220 844 4230
rect 1012 4144 1112 4154
rect 1012 3982 1112 4044
rect 1202 4144 1302 4407
rect 1202 4034 1302 4044
rect 1470 4330 1570 4340
rect 1470 3982 1570 4230
rect 1660 4144 1760 4407
rect 1660 4034 1760 4044
rect 1928 4330 2028 4340
rect 1928 3982 2028 4230
rect 2118 4330 2218 4407
rect 2118 4220 2218 4230
rect 2386 4144 2486 4154
rect 2386 3982 2486 4044
rect 912 3972 1112 3982
rect 912 3910 1112 3920
rect 1370 3972 1570 3982
rect 1370 3910 1570 3920
rect 1828 3972 2028 3982
rect 1828 3910 2028 3920
rect 2286 3972 2486 3982
rect 2286 3910 2486 3920
rect 650 3869 744 3879
rect 650 3722 744 3732
rect 2485 3869 2579 3879
rect 2485 3722 2579 3732
rect 557 3667 615 3677
rect 1569 3611 1663 3621
rect 1131 3463 1183 3473
rect 1569 3464 1663 3474
rect 2047 3463 2099 3473
rect 1183 3303 2047 3394
rect 2879 3394 2979 4993
rect 3048 4876 4426 4886
rect 3861 4602 3913 4876
rect 3861 4521 3913 4531
rect 4217 4602 4269 4876
rect 4217 4521 4269 4531
rect 4305 4497 4357 4507
rect 3949 4382 4001 4392
rect 2099 3303 2979 3394
rect 1131 3294 2979 3303
rect 3644 4052 3748 4062
rect 1131 3293 1183 3294
rect 2047 3293 2099 3294
rect 615 3129 2685 3139
rect 557 3016 2685 3026
rect -766 2896 3644 2903
rect -801 2893 3644 2896
rect 3949 3917 4001 4303
rect 3949 3707 4001 3717
rect 4305 4253 4357 4426
rect 4588 4253 4660 5369
rect 4305 4181 4779 4253
rect 4305 3917 4357 4181
rect 4305 3707 4357 3717
rect 3821 3621 3873 3631
rect 3748 3421 3821 3553
rect 4177 3621 4229 3631
rect 3873 3421 4177 3553
rect 3748 3411 4229 3421
rect -801 2886 -766 2893
rect -863 594 -801 604
rect -684 2786 3748 2796
rect 546 2494 598 2786
rect -518 2218 -454 2228
rect 1598 2494 1662 2504
rect 1598 2284 1662 2294
rect 2662 2494 2714 2786
rect 546 2184 598 2194
rect 2662 2184 2714 2194
rect 3714 2218 3778 2228
rect -518 2008 -454 2018
rect 3714 2008 3778 2018
rect -441 1968 199 1978
rect -441 1906 199 1916
rect 617 1968 1257 1978
rect 617 1906 1257 1916
rect 1675 1968 2315 1978
rect 1675 1906 2315 1916
rect 2733 1968 3373 1978
rect 2733 1906 3373 1916
rect -441 1812 -341 1906
rect -441 1702 -341 1712
rect 427 1630 527 1640
rect 427 1444 527 1530
rect 617 1630 717 1906
rect 617 1520 717 1530
rect 1485 1812 1585 1822
rect 1485 1444 1585 1712
rect 1675 1630 1775 1906
rect 1675 1520 1775 1530
rect 2543 1812 2643 1822
rect -113 1434 527 1444
rect -113 1372 527 1382
rect 945 1434 1585 1444
rect 2543 1443 2643 1712
rect 2733 1812 2833 1906
rect 2733 1702 2833 1712
rect 3601 1630 3701 1640
rect 3601 1444 3701 1530
rect 945 1372 1585 1382
rect 2003 1433 2643 1443
rect 2003 1371 2643 1381
rect 3061 1434 3701 1444
rect 3061 1372 3701 1382
rect 3983 1407 4080 1417
rect -518 1332 -454 1342
rect 3714 1332 3778 1342
rect -518 1122 -454 1132
rect 546 1156 598 1166
rect 2662 1156 2714 1166
rect 546 604 598 856
rect 1598 1056 1662 1066
rect 1598 846 1662 856
rect 3714 1122 3778 1132
rect 2662 604 2714 856
rect -684 603 3941 604
rect -684 594 3983 603
rect 3941 593 3983 594
rect 4080 602 4099 603
rect 4080 593 4217 602
rect -863 228 3840 229
rect 4099 228 4217 593
rect -863 219 4217 228
rect 3840 218 4217 219
rect 4079 217 4217 218
<< via2 >>
rect 1008 5713 1064 5853
rect 3138 5368 3279 5430
rect 1568 4732 1662 4869
rect 651 4521 745 4658
rect 2483 4521 2577 4658
rect 650 3732 744 3869
rect 2485 3732 2579 3869
rect 1569 3474 1663 3611
rect -518 2018 -454 2218
rect 1598 2294 1662 2494
rect 3714 2018 3778 2218
rect -518 1132 -454 1332
rect 1598 856 1662 1056
rect 3714 1132 3778 1332
<< metal3 >>
rect 2618 6927 2867 7034
rect 998 5853 1074 5858
rect 998 5768 1008 5853
rect 220 5713 1008 5768
rect 1064 5713 1074 5853
rect 220 5708 1074 5713
rect 3128 5433 3289 5435
rect 3128 5365 3138 5433
rect 3279 5365 3289 5433
rect 3128 5363 3289 5365
rect 1558 4869 2905 4874
rect 1558 4732 1568 4869
rect 1662 4732 2905 4869
rect 1558 4727 1672 4732
rect 641 4658 755 4663
rect 641 4521 651 4658
rect 745 4521 755 4658
rect 641 4516 755 4521
rect 2473 4658 2587 4663
rect 2473 4521 2483 4658
rect 2577 4521 2587 4658
rect 2473 4516 2587 4521
rect 2758 3874 2905 4732
rect 640 3869 2905 3874
rect 640 3732 650 3869
rect 744 3732 2485 3869
rect 2579 3732 2905 3869
rect 640 3727 2905 3732
rect 1559 3611 1673 3616
rect 1559 3474 1569 3611
rect 1663 3474 1673 3611
rect 1559 3469 1673 3474
rect 2758 2499 2905 3727
rect 1588 2494 4228 2499
rect 1588 2294 1598 2494
rect 1662 2399 4228 2494
rect 1662 2294 1672 2399
rect 1588 2289 1672 2294
rect -528 2218 -444 2223
rect -528 2018 -518 2218
rect -454 2018 -444 2218
rect -528 2013 -444 2018
rect 3704 2218 3788 2223
rect 3704 2018 3714 2218
rect 3778 2018 3788 2218
rect 3704 2013 3788 2018
rect 4128 1337 4228 2399
rect -528 1332 4228 1337
rect -528 1132 -518 1332
rect -454 1237 3714 1332
rect -454 1132 -444 1237
rect -528 1127 -444 1132
rect 3704 1132 3714 1237
rect 3778 1237 4228 1332
rect 3778 1132 3788 1237
rect 3704 1127 3788 1132
rect 1588 1056 1672 1061
rect 1588 856 1598 1056
rect 1662 856 1672 1056
rect 1588 851 1672 856
<< via3 >>
rect 3138 5430 3279 5433
rect 3138 5368 3279 5430
rect 3138 5365 3279 5368
rect 651 4521 745 4658
rect 2483 4521 2577 4658
rect 1569 3474 1663 3611
rect -518 2018 -454 2218
rect 3714 2018 3778 2218
rect 1598 856 1662 1056
<< metal4 >>
rect 3129 5434 3240 6046
rect 3129 5433 3280 5434
rect 3129 5365 3138 5433
rect 3279 5430 3280 5433
rect 3279 5368 3348 5430
rect 3279 5365 3280 5368
rect 3129 5364 3280 5365
rect 374 4658 2578 4659
rect 374 4521 651 4658
rect 745 4521 2483 4658
rect 2577 4521 2578 4658
rect 374 4520 2578 4521
rect 374 3612 513 4520
rect 374 3611 1686 3612
rect 374 3474 1569 3611
rect 1663 3474 1686 3611
rect 374 3473 1686 3474
rect -519 2218 -453 2219
rect -519 2117 -518 2218
rect -971 2018 -518 2117
rect -454 2117 -453 2218
rect 374 2117 513 3473
rect 3713 2218 3779 2219
rect 3713 2117 3714 2218
rect -454 2018 3714 2117
rect 3778 2018 3779 2218
rect -971 2017 3779 2018
rect -971 955 -871 2017
rect 1597 1056 1663 1057
rect 1597 955 1598 1056
rect -971 856 1598 955
rect 1662 856 1663 1056
rect -971 855 1663 856
use sky130_fd_pr__nfet_01v8_lvt_D5AAWA  sky130_fd_pr__nfet_01v8_lvt_D5AAWA_0
timestamp 1741119366
transform 1 0 2302 0 1 4798
box -258 -388 258 388
use sky130_fd_pr__nfet_01v8_lvt_RX9YJP  sky130_fd_pr__nfet_01v8_lvt_RX9YJP_0
timestamp 1741136105
transform 1 0 4287 0 1 4514
box -73 -188 73 188
use sky130_fd_pr__pfet_01v8_lvt_227YHS  sky130_fd_pr__pfet_01v8_lvt_227YHS_0
timestamp 1741123092
transform 1 0 3217 0 1 1094
box -594 -350 594 350
use sky130_fd_pr__cap_mim_m3_1_Q3FE5R  XC2
timestamp 1741058913
transform 1 0 4726 0 1 7694
box -1886 -1740 1886 1740
use sky130_fd_pr__nfet_01v8_lvt_D5AAWA  XM1
timestamp 1741119366
transform 1 0 928 0 1 4798
box -258 -388 258 388
use sky130_fd_pr__nfet_01v8_lvt_D5AAWA  XM2
timestamp 1741119366
transform 1 0 928 0 1 3591
box -258 -388 258 388
use sky130_fd_pr__nfet_01v8_22NDE3  XM3
timestamp 1741058913
transform 0 -1 1641 1 0 6011
box -525 -760 525 760
use sky130_fd_pr__pfet_01v8_lvt_227YHS  XM4
timestamp 1741123092
transform 1 0 43 0 1 2256
box -594 -350 594 350
use sky130_fd_pr__pfet_01v8_lvt_227YHS  XM5
timestamp 1741123092
transform 1 0 43 0 1 1094
box -594 -350 594 350
use sky130_fd_pr__pfet_01v8_lvt_K7KF7V  XM6
timestamp 1741058913
transform 1 0 4267 0 1 3669
box -231 -479 231 479
use sky130_fd_pr__pfet_01v8_lvt_K7KF7V  XM7
timestamp 1741058913
transform 1 0 3911 0 1 3669
box -231 -479 231 479
use sky130_fd_pr__nfet_01v8_lvt_RX9YJP  XM9
timestamp 1741136105
transform 1 0 3931 0 1 4514
box -73 -188 73 188
use sky130_fd_pr__pfet_01v8_lvt_227YHS  XM10
timestamp 1741123092
transform 1 0 1101 0 1 2256
box -594 -350 594 350
use sky130_fd_pr__pfet_01v8_lvt_227YHS  XM11
timestamp 1741123092
transform 1 0 2159 0 1 2256
box -594 -350 594 350
use sky130_fd_pr__pfet_01v8_lvt_227YHS  XM13
timestamp 1741123092
transform 1 0 1101 0 1 1094
box -594 -350 594 350
use sky130_fd_pr__pfet_01v8_lvt_227YHS  XM14
timestamp 1741123092
transform 1 0 2159 0 1 1094
box -594 -350 594 350
use sky130_fd_pr__pfet_01v8_lvt_227YHS  XM15
timestamp 1741123092
transform 1 0 3217 0 1 2256
box -594 -350 594 350
use sky130_fd_pr__nfet_01v8_lvt_D5AAWA  XM16
timestamp 1741119366
transform 1 0 1386 0 1 4798
box -258 -388 258 388
use sky130_fd_pr__nfet_01v8_lvt_D5AAWA  XM17
timestamp 1741119366
transform 1 0 1844 0 1 4798
box -258 -388 258 388
use sky130_fd_pr__nfet_01v8_lvt_D5AAWA  XM18
timestamp 1741119366
transform 1 0 2302 0 1 3591
box -258 -388 258 388
use sky130_fd_pr__nfet_01v8_lvt_D5AAWA  XM19
timestamp 1741119366
transform 1 0 1386 0 1 3591
box -258 -388 258 388
use sky130_fd_pr__nfet_01v8_lvt_D5AAWA  XM20
timestamp 1741119366
transform 1 0 1844 0 1 3591
box -258 -388 258 388
use sky130_fd_pr__res_xhigh_po_0p35_NX66A7  XR1
timestamp 1741058913
transform 0 -1 3862 1 0 5405
box -201 -702 201 702
<< labels >>
rlabel metal2 4215 390 4215 390 3 vcc
port 1 e
rlabel metal2 463 6644 463 6644 7 vss
port 2 w
rlabel metal2 4778 4214 4778 4214 3 vo3
port 3 e
rlabel metal1 -66 4276 -66 4276 7 vd3
port 4 w
rlabel metal1 -66 4099 -66 4099 7 vd4
port 5 w
rlabel metal3 2619 6975 2619 6975 7 vd1
port 7 w
rlabel metal3 221 5737 221 5737 7 vb
port 6 w
<< end >>
