** sch_path: /home/zerotoasic/Dalin/Projects/tinytape/voltage_ref_BJT/BGR_BJT_final.sch
.subckt BGR_BJT_final vcc vref vss
*.PININFO vcc:I vss:I vref:O
x1 vcc net1 net2 vss BGR_BJT_stage1
x2 vcc net1 vref net2 vss BGR_BJT_stage2
.ends

* expanding   symbol:  /home/zerotoasic/Dalin/Projects/tinytape/voltage_ref_BJT/BGR_BJT_stage1.sym # of pins=4
** sym_path: /home/zerotoasic/Dalin/Projects/tinytape/voltage_ref_BJT/BGR_BJT_stage1.sym
** sch_path: /home/zerotoasic/Dalin/Projects/tinytape/voltage_ref_BJT/BGR_BJT_stage1.sch
.subckt BGR_BJT_stage1 vcc vr vref0 vss
*.PININFO vcc:I vref0:O vr:O vss:I
XM1 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM2 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM3 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM8 vr vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 m=1
XM9 net2 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM4 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM5 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM6 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM7 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM10 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM11 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM12 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM14 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM15 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM16 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM17 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM18 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM19 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM20 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM21 vr net2 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM22 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM23 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM24 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM25 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM26 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM27 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM28 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM29 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM30 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM31 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM32 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM33 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM34 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM35 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM36 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM37 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM38 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM39 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM40 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM41 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM42 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM43 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM44 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM45 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM46 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM47 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM48 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM49 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM50 vref0 net2 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM51 net1 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM52 vr vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 m=1
XQ1 vss vss net2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XM13 net2 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  /home/zerotoasic/Dalin/Projects/tinytape/voltage_ref_BJT/BGR_BJT_stage2.sym # of pins=5
** sym_path: /home/zerotoasic/Dalin/Projects/tinytape/voltage_ref_BJT/BGR_BJT_stage2.sym
** sch_path: /home/zerotoasic/Dalin/Projects/tinytape/voltage_ref_BJT/BGR_BJT_stage2.sch
.subckt BGR_BJT_stage2 vcc vr vref vref0 vss
*.PININFO vref:O vcc:I vss:I vref0:I vr:I
XM4 net2 net3 vref0 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM5 net3 net3 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM6 net1 net4 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM7 net4 net4 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM10 net3 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM11 net4 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM12 vref vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM16 net5 net6 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM15 net6 net6 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM14 net6 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM19 vref net7 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM18 net7 net7 vref vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM17 net7 vr vcc vcc sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 m=1
XM1 net3 net3 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM2 net3 net3 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM3 net3 net3 net2 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM8 net4 net4 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM9 net4 net4 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM13 net4 net4 net1 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM20 net6 net6 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM21 net6 net6 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM22 net6 net6 net5 vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM23 net7 net7 vref vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM24 net7 net7 vref vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM25 net7 net7 vref vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
.ends

.end
