* NGSPICE file created from 3_OTA_flat.ext - technology: sky130A

.subckt x3_OTA_flat vo3 vin_p vin_n vcc vss
X0 a_9040_n3397# 3rd_3_OTA_0.vd3.t12 a_7434_495.t3 vss.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=34800,1316 d=17400,658
X1 a_n1236_n9479.t47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X2 a_7434_1657.t3 3rd_3_OTA_0.vd4.t8 a_9040_n3397# vss.t36 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=17400,658
X3 3rd_3_OTA_0.vd3.t11 OTA_stage1_0.vd2.t3 a_n1050_166.t5 vcc.t29 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X4 OTA_stage1_0.vd2.t0 vin_p.t0 a_n10077_1624# vss.t61 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X5 vo3.t1 a_7434_1657.t12 vcc.t20 vcc.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.6 l=0.35
**devattr s=30160,1156 d=30160,1156
X6 a_n1236_n9479.t46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X7 a_n1236_n9479.t45 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X8 a_7434_1657.t9 a_7434_1657.t8 vcc.t18 vcc.t17 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X9 a_7434_495.t11 a_7434_495.t10 vcc.t47 vcc.t15 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=29000,1116
X10 OTA_vref_0.vb1.t4 a_2382_n6868# a_2470_n7958# vss.t13 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X11 a_n1236_n9479.t44 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X12 a_2382_n8158# OTA_vref_0.OTA_vref_stage2_0.vr.t20 vcc.t49 vcc.t48 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X13 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 a_n1236_n9479.t43 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X14 a_11847_n1701# a_11847_n1701# vss.t23 vss.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X15 vss.t37 3rd_3_OTA_0.vd3.t5 3rd_3_OTA_0.vd3.t6 vss.t26 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X16 a_11275_n2439.t1 3rd_3_OTA_0.vd1 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X17 OTA_stage1_0.vd2.t2 OTA_stage1_0.vd2.t0 vcc.t28 vcc.t26 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X18 vss.t43 a_n1236_n9479.t30 a_n1236_n9479.t31 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X19 3rd_3_OTA_0.vb a_2382_n4288# a_2382_n4288# vss.t51 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X20 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 a_n1236_n9479.t42 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X21 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 a_n1236_n9479.t41 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X22 vss.t0 vss.t14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X23 3rd_3_OTA_0.vd1.t1 OTA_stage1_0.vd2.t0 vcc.t27 vcc.t26 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X24 a_n10077_1624# vin_p.t1 OTA_stage1_0.vd2.t0 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X25 a_7434_1657.t7 a_7434_1657.t6 vcc.t16 vcc.t15 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=29000,1116
X26 vss.t59 a_n1236_n9479.t28 a_n1236_n9479.t29 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X27 a_11847_n1701# a_7434_495.t12 vcc.t46 vcc.t45 sky130_fd_pr__pfet_01v8_lvt ad=0.754 pd=5.78 as=0 ps=0 w=2.6 l=0.35
**devattr s=30160,1156 d=30160,1156
X28 a_7434_495.t2 3rd_3_OTA_0.vd3.t13 a_9040_n3397# vss.t36 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=17400,658
X29 a_2382_n6868# a_2382_n6868# OTA_vref_0.vb1.t3 vss.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X30 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 a_n1236_n9479.t40 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X31 OTA_vref_0.OTA_vref_stage2_0.vr.t19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X32 3rd_3_OTA_0.vd3.t8 3rd_3_OTA_0.vd3.t7 vss.t35 vss.t30 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X33 vcc.t14 a_7434_1657.t10 a_7434_1657.t11 vcc.t13 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X34 a_2470_n7958# a_2382_n8158# a_2382_n8158# vss.t56 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X35 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 a_n1236_n9479.t39 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X36 OTA_vref_0.OTA_vref_stage2_0.vr.t18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X37 a_n1050_166.t4 OTA_stage1_0.vd2.t4 3rd_3_OTA_0.vd3.t10 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X38 a_2382_n6868# a_2382_n6868# OTA_vref_0.vb1.t2 vss.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X39 vcc.t12 a_7434_1657.t4 a_7434_1657.t5 vcc.t11 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=29000,1116 d=14500,558
X40 a_2382_n4288# a_2382_n4288# 3rd_3_OTA_0.vb vss.t50 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=5800,258 d=5800,258
X41 a_n1236_n9479.t38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X42 a_n1050_166.t10 OTA_vref_0.vb1.t6 vcc.t41 vcc.t40 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=81200,2916
X43 3rd_3_OTA_0.vd4.t9 3rd_3_OTA_0.vd1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X44 vss.t62 a_n1236_n9479.t26 a_n1236_n9479.t27 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X45 OTA_vref_0.OTA_vref_stage2_0.vr.t17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X46 OTA_vref_0.OTA_vref_stage2_0.vr.t16 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X47 OTA_vref_0.OTA_vref_stage2_0.vr.t3 OTA_vref_0.OTA_vref_stage2_0.vr.t2 vcc.t34 vcc.t9 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=2900,158 d=5800,316
X48 vss.t34 3rd_3_OTA_0.vd3.t14 3rd_3_OTA_0.vd4.t4 vss.t28 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X49 OTA_vref_0.vb1.t1 a_2382_n6868# a_2382_n6868# vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X50 vcc.t36 OTA_vref_0.vb1.t7 a_n1050_166.t8 vcc.t35 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X51 vss.t8 a_n1236_n9479.t24 a_n1236_n9479.t25 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X52 a_9040_n3397# 3rd_3_OTA_0.vd4.t10 a_7434_1657.t2 vss.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=34800,1316 d=17400,658
X53 3rd_3_OTA_0.vb a_2382_n4288# a_2470_n5378# vss.t49 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X54 a_2382_n5578# OTA_vref_0.OTA_vref_stage2_0.vr.t21 vcc.t8 vcc.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X55 vss.t46 a_n1236_n9479.t22 a_n1236_n9479.t23 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X56 vss.t44 a_n1236_n9479.t20 a_n1236_n9479.t21 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X57 a_n1050_166.t1 3rd_3_OTA_0.vd1.t4 3rd_3_OTA_0.vd4.t0 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X58 vss.t60 a_n1236_n9479.t18 a_n1236_n9479.t19 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X59 a_n10077_1624# vin_n.t0 3rd_3_OTA_0.vd1.t3 vss.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X60 a_2470_n7958# a_2382_n8158# OTA_vref_0.OTA_vref_stage2_0.vref0.t32 vss.t55 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X61 vcc.t39 OTA_vref_0.vb1.t8 a_n1050_166.t9 vcc.t38 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=81200,2916 d=40600,1458
X62 a_n1050_166.t6 3rd_3_OTA_0.vd1.t5 3rd_3_OTA_0.vd4.t5 vcc.t25 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X63 3rd_3_OTA_0.vd3.t2 3rd_3_OTA_0.vd3.t1 vss.t33 vss.t26 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X64 a_n1236_n9479.t17 a_n1236_n9479.t16 vss.t4 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X65 a_2382_n4288# a_2382_n4288# 3rd_3_OTA_0.vb vss.t48 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=5800,258 d=5800,258
X66 OTA_vref_0.OTA_vref_stage2_0.vr.t15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X67 vss.t7 a_n1236_n9479.t14 a_n1236_n9479.t15 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X68 a_n1050_166.t3 OTA_stage1_0.vd2.t5 3rd_3_OTA_0.vd3.t0 vcc.t25 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X69 a_n1236_n9479.t13 a_n1236_n9479.t12 vss.t2 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X70 a_2470_n5378# a_2382_n5578# a_2382_n5578# vss.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X71 vcc.t6 OTA_vref_0.OTA_vref_stage2_0.vr.t22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 vcc.t5 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X72 vss.t32 3rd_3_OTA_0.vd3.t15 3rd_3_OTA_0.vd4.t3 vss.t26 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X73 OTA_vref_0.OTA_vref_stage2_0.vr.t14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X74 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 OTA_vref_0.OTA_vref_stage2_0.vr.t13 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X75 OTA_vref_0.OTA_vref_stage2_0.vr.t12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X76 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 OTA_vref_0.OTA_vref_stage2_0.vr.t11 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X77 a_7434_1657.t1 3rd_3_OTA_0.vd4.t11 a_9040_n3397# vss.t24 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=34800,1316
X78 3rd_3_OTA_0.vd3.t9 OTA_stage1_0.vd2.t6 a_n1050_166.t2 vcc.t24 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X79 a_2382_n8158# a_2382_n8158# a_2470_n7958# vss.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X80 3rd_3_OTA_0.vd1.t2 vin_n.t1 a_n10077_1624# vss.t41 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X81 a_2382_n5578# a_2382_n5578# a_2470_n5378# vss.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X82 a_7434_495.t9 a_7434_495.t8 vcc.t44 vcc.t17 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X83 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 a_n1236_n9479.t37 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X84 3rd_3_OTA_0.vb a_2382_n4288# a_2382_n4288# vss.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=11600,516
X85 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 OTA_vref_0.OTA_vref_stage2_0.vr.t10 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X86 a_n1050_166.t0 OTA_vref_0.vb1.t9 vcc.t3 vcc.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 OTA_vref_0.OTA_vref_stage2_0.vr.t23 vcc.t33 vcc.t32 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=11600,516
X88 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 OTA_vref_0.OTA_vref_stage2_0.vr.t9 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X89 a_2470_n5378# a_2382_n5578# OTA_vref_0.vb1.t5 vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X90 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 OTA_vref_0.OTA_vref_stage2_0.vr.t8 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X91 a_2382_n6868# OTA_vref_0.OTA_vref_stage2_0.vr.t24 vcc.t31 vcc.t30 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X92 a_n1236_n9479.t11 a_n1236_n9479.t10 vss.t3 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X93 a_2470_n7958# a_2382_n8158# a_2382_n8158# vss.t53 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X94 vcc.t43 a_7434_495.t4 a_7434_495.t5 vcc.t13 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=14500,558 d=14500,558
X95 3rd_3_OTA_0.vd4.t2 3rd_3_OTA_0.vd3.t16 vss.t31 vss.t30 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X96 a_n1236_n9479.t9 a_n1236_n9479.t8 vss.t57 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X97 a_n1236_n9479.t7 a_n1236_n9479.t6 vss.t45 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X98 vo3.t2 a_11847_n1701# vss.t21 vss.t20 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X99 a_9040_n3397# 3rd_3_OTA_0.vd4.t12 a_7434_1657.t0 vss.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=17400,658 d=17400,658
X100 vss.t29 3rd_3_OTA_0.vd3.t3 3rd_3_OTA_0.vd3.t4 vss.t28 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X101 a_2382_n8158# a_2382_n8158# a_2470_n7958# vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X102 a_n1236_n9479.t5 a_n1236_n9479.t4 vss.t42 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X103 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 OTA_vref_0.OTA_vref_stage2_0.vr.t7 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X104 vcc.t23 OTA_stage1_0.vd2.t0 3rd_3_OTA_0.vd1.t0 vcc.t21 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X105 vcc.t10 OTA_vref_0.OTA_vref_stage2_0.vr.t0 OTA_vref_0.OTA_vref_stage2_0.vr.t1 vcc.t9 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=5800,316 d=2900,158
X106 a_n1236_n9479.t36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X107 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 a_n1236_n9479.t35 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X108 a_2382_n5578# a_2382_n5578# a_2470_n5378# vss.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X109 a_n1236_n9479.t3 a_n1236_n9479.t2 vss.t40 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X110 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 a_n1236_n9479.t34 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X111 3rd_3_OTA_0.vd4.t7 3rd_3_OTA_0.vd1.t6 a_n1050_166.t11 vcc.t24 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X112 OTA_vref_0.vb1.t0 a_2382_n6868# a_2382_n6868# vss.t9 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X113 3rd_3_OTA_0.vb OTA_vref_0.OTA_vref_stage2_0.vr.t25 vcc.t1 vcc.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X114 3rd_3_OTA_0.vd4.t6 3rd_3_OTA_0.vd1.t7 a_n1050_166.t7 vcc.t29 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X115 vcc.t22 OTA_stage1_0.vd2.t0 OTA_stage1_0.vd2.t1 vcc.t21 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X116 vcc.t42 a_7434_495.t6 a_7434_495.t7 vcc.t11 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.5 l=5
**devattr s=29000,1116 d=14500,558
X117 a_9040_n3397# 3rd_3_OTA_0.vb vss.t67 vss.t63 sky130_fd_pr__nfet_01v8 ad=1.048143 pd=7.775429 as=0 ps=0 w=5.5 l=1.5
**devattr s=31900,1158 d=63800,2316
X118 OTA_vref_0.OTA_vref_stage2_0.vref0.t0 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 OTA_vref_0.OTA_vref_stage2_0.vr.t6 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X119 3rd_3_OTA_0.vd4.t1 3rd_3_OTA_0.vd3.t17 vss.t27 vss.t26 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X120 a_n1236_n9479.t33 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X121 a_n10077_1624# 3rd_3_OTA_0.vb vss.t66 vss.t65 sky130_fd_pr__nfet_01v8 ad=0.483333 pd=3.526667 as=0 ps=0 w=3 l=5
**devattr s=34800,1316 d=34800,1316
X122 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 OTA_vref_0.OTA_vref_stage2_0.vr.t5 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X123 a_9040_n3397# 3rd_3_OTA_0.vd3.t18 a_7434_495.t1 vss.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.571714 pd=4.241143 as=0 ps=0 w=3 l=2
**devattr s=17400,658 d=17400,658
X124 a_n1236_n9479.t32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X125 a_11275_n2439.t0 vo3.t0 vss.t5 sky130_fd_pr__res_xhigh_po_0p35 l=1.2
X126 a_2382_n4288# OTA_vref_0.OTA_vref_stage2_0.vr.t26 vcc.t37 vcc.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=2
**devattr s=11600,516 d=11600,516
X127 OTA_vref_0.OTA_vref_stage2_0.vr.t4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X128 a_7434_495.t0 3rd_3_OTA_0.vd3.t19 a_9040_n3397# vss.t24 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.571714 ps=4.241143 w=3 l=2
**devattr s=17400,658 d=34800,1316
X129 vss.t64 3rd_3_OTA_0.vb a_9040_n3397# vss.t63 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=1.048143 ps=7.775429 w=5.5 l=1.5
**devattr s=63800,2316 d=31900,1158
X130 a_2470_n5378# a_2382_n5578# a_2382_n5578# vss.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X131 a_n1236_n9479.t1 a_n1236_n9479.t0 vss.t39 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
R0 3rd_3_OTA_0.vd3.n2 3rd_3_OTA_0.vd3.t8 60.3532
R1 3rd_3_OTA_0.vd3.n1 3rd_3_OTA_0.vd3.t4 60.3532
R2 3rd_3_OTA_0.vd3.n3 3rd_3_OTA_0.vd3.n10 48.5755
R3 3rd_3_OTA_0.vd3.n0 3rd_3_OTA_0.vd3.t19 44.0616
R4 3rd_3_OTA_0.vd3.n0 3rd_3_OTA_0.vd3.t13 44.0379
R5 3rd_3_OTA_0.vd3.n0 3rd_3_OTA_0.vd3.t18 44.0379
R6 3rd_3_OTA_0.vd3 3rd_3_OTA_0.vd3.t12 43.8241
R7 3rd_3_OTA_0.vd3.n5 3rd_3_OTA_0.vd3.t0 19.1315
R8 3rd_3_OTA_0.vd3.n5 3rd_3_OTA_0.vd3.t11 18.308
R9 3rd_3_OTA_0.vd3.n5 3rd_3_OTA_0.vd3.n6 16.2734
R10 3rd_3_OTA_0.vd3.n13 3rd_3_OTA_0.vd3.n1 14.6534
R11 3rd_3_OTA_0.vd3.n10 3rd_3_OTA_0.vd3.t6 11.6005
R12 3rd_3_OTA_0.vd3.n10 3rd_3_OTA_0.vd3.t2 11.6005
R13 3rd_3_OTA_0.vd3 3rd_3_OTA_0.vd3.n1 11.2227
R14 3rd_3_OTA_0.vd3.n3 3rd_3_OTA_0.vd3.n7 8.08817
R15 3rd_3_OTA_0.vd3 3rd_3_OTA_0.vd3.n2 7.9105
R16 3rd_3_OTA_0.vd3.n8 3rd_3_OTA_0.vd3.t7 3.58326
R17 3rd_3_OTA_0.vd3.n9 3rd_3_OTA_0.vd3.t15 3.58326
R18 3rd_3_OTA_0.vd3.n11 3rd_3_OTA_0.vd3.t17 3.58326
R19 3rd_3_OTA_0.vd3.n12 3rd_3_OTA_0.vd3.t3 3.58326
R20 3rd_3_OTA_0.vd3.n8 3rd_3_OTA_0.vd3.t16 3.58267
R21 3rd_3_OTA_0.vd3.n9 3rd_3_OTA_0.vd3.t5 3.58267
R22 3rd_3_OTA_0.vd3.n11 3rd_3_OTA_0.vd3.t1 3.58267
R23 3rd_3_OTA_0.vd3.n12 3rd_3_OTA_0.vd3.t14 3.58267
R24 3rd_3_OTA_0.vd3.n4 3rd_3_OTA_0.vd3.n13 3.54985
R25 3rd_3_OTA_0.vd3.n7 3rd_3_OTA_0.vd3.n5 2.67636
R26 3rd_3_OTA_0.vd3.n1 3rd_3_OTA_0.vd3.n12 2.60735
R27 3rd_3_OTA_0.vd3.n2 3rd_3_OTA_0.vd3.n8 2.58162
R28 3rd_3_OTA_0.vd3 3rd_3_OTA_0.vd3.n0 2.5555
R29 3rd_3_OTA_0.vd3 3rd_3_OTA_0.vd3.n7 2.29713
R30 3rd_3_OTA_0.vd3.n6 3rd_3_OTA_0.vd3.t10 1.90483
R31 3rd_3_OTA_0.vd3.n6 3rd_3_OTA_0.vd3.t9 1.90483
R32 3rd_3_OTA_0.vd3.n2 3rd_3_OTA_0.vd3.n4 1.69798
R33 3rd_3_OTA_0.vd3.n13 3rd_3_OTA_0.vd3.n11 1.61224
R34 3rd_3_OTA_0.vd3.n4 3rd_3_OTA_0.vd3.n9 1.61224
R35 3rd_3_OTA_0.vd3.n4 3rd_3_OTA_0.vd3.n3 1.22519
R36 a_7434_495.n1 a_7434_495.t12 387.724
R37 a_7434_495.n13 a_7434_495.t11 96.4663
R38 a_7434_495.n10 a_7434_495.n9 84.9005
R39 a_7434_495.n17 a_7434_495.t0 38.5275
R40 a_7434_495.t3 a_7434_495.n17 37.908
R41 a_7434_495.n16 a_7434_495.n15 32.1023
R42 a_7434_495.n8 a_7434_495.t8 13.386
R43 a_7434_495.n7 a_7434_495.t4 13.3552
R44 a_7434_495.n12 a_7434_495.t10 13.3552
R45 a_7434_495.n4 a_7434_495.t6 13.3139
R46 a_7434_495.n9 a_7434_495.t5 11.4265
R47 a_7434_495.n9 a_7434_495.t9 11.4265
R48 a_7434_495.n0 a_7434_495.n4 7.96494
R49 a_7434_495.n11 a_7434_495.n2 6.81377
R50 a_7434_495.n14 a_7434_495.n13 6.51669
R51 a_7434_495.n1 a_7434_495.n7 5.8066
R52 a_7434_495.n15 a_7434_495.t1 5.8005
R53 a_7434_495.n15 a_7434_495.t2 5.8005
R54 a_7434_495.n8 a_7434_495.n0 5.77549
R55 a_7434_495.n12 a_7434_495.n1 5.58783
R56 a_7434_495.n4 a_7434_495.n3 0.495597
R57 a_7434_495.n3 a_7434_495.n2 4.99728
R58 a_7434_495.n10 a_7434_495.n5 0.783109
R59 a_7434_495.n7 a_7434_495.n5 0.638655
R60 a_7434_495.n7 a_7434_495.n6 0.592891
R61 a_7434_495.n6 a_7434_495.n8 0.541261
R62 a_7434_495.n8 a_7434_495.n5 0.510015
R63 a_7434_495.n13 a_7434_495.n12 0.501908
R64 a_7434_495.n16 a_7434_495.n14 0.47591
R65 a_7434_495.n14 a_7434_495.n2 0.4047
R66 a_7434_495.n17 a_7434_495.n16 0.393745
R67 a_7434_495.n6 a_7434_495.n11 0.293331
R68 a_7434_495.n11 a_7434_495.n10 0.25257
R69 a_7434_495.t7 a_7434_495.n3 96.4689
R70 a_7434_495.n1 a_7434_495.n0 1.5605
R71 vss.n53 vss.t26 6.51798e+06
R72 vss.n311 vss.n57 5.4843e+06
R73 vss.n57 vss.n54 3.3e+06
R74 vss.n54 vss.n53 2.376e+06
R75 vss.n313 vss.n312 1.23016e+06
R76 vss.n313 vss.n54 402600
R77 vss.n312 vss.n311 354428
R78 vss.n367 vss.n315 156933
R79 vss.n465 vss.n6 147329
R80 vss.n336 vss.n315 114006
R81 vss.n466 vss.n465 72897.2
R82 vss.t26 vss.n6 36497.6
R83 vss.n467 vss.n466 31912.6
R84 vss.n463 vss.n7 27614.8
R85 vss.n463 vss.n8 27609
R86 vss.n450 vss.n7 27609
R87 vss.n450 vss.n8 27603.2
R88 vss.n443 vss.n33 26954.2
R89 vss.n422 vss.n33 26954.2
R90 vss.n443 vss.n34 26948.4
R91 vss.n422 vss.n34 26948.4
R92 vss.n437 vss.n424 25442
R93 vss.n424 vss.n423 25442
R94 vss.n437 vss.n425 25436.2
R95 vss.n425 vss.n423 25436.2
R96 vss.n336 vss.n6 24232.3
R97 vss.n447 vss.n28 17753.2
R98 vss.n447 vss.n29 17753.2
R99 vss.n309 vss.n28 17753.2
R100 vss.n309 vss.n29 17753.2
R101 vss.n466 vss.n5 16119.1
R102 vss.n317 vss.n316 12277.7
R103 vss.n398 vss.n316 12277.7
R104 vss.n397 vss.n317 12277.7
R105 vss.n398 vss.n397 12277.7
R106 vss.n337 vss.n336 9391.71
R107 vss.n394 vss.n49 6732.77
R108 vss.n401 vss.n49 6732.77
R109 vss.n394 vss.n50 6732.77
R110 vss.n401 vss.n50 6732.77
R111 vss.n367 vss.n337 6373.53
R112 vss.n432 vss.n3 6275.03
R113 vss.n468 vss.n3 6275.03
R114 vss.n432 vss.n4 6275.03
R115 vss.n468 vss.n4 6275.03
R116 vss.n57 vss.n56 5636.95
R117 vss.n53 vss.n52 5636.95
R118 vss.n347 vss.n334 4519.41
R119 vss.n347 vss.n335 4519.41
R120 vss.n369 vss.n334 4519.41
R121 vss.n369 vss.n335 4519.41
R122 vss.n465 vss.n464 4064.84
R123 vss.n344 vss.n338 3412.74
R124 vss.n344 vss.n339 3412.74
R125 vss.n365 vss.n338 3406.94
R126 vss.n365 vss.n339 3406.94
R127 vss.n346 vss.n337 2223.62
R128 vss.n449 vss.n448 2022.67
R129 vss.n372 vss.n332 1960.4
R130 vss.n440 vss.n439 1944.26
R131 vss.t41 vss.n5 1579.6
R132 vss.n430 vss.t58 1579.6
R133 vss.n220 vss.t0 1564.71
R134 vss.n439 vss.t61 1324.96
R135 vss.n438 vss.t6 1324.96
R136 vss.n261 vss.n94 1305.6
R137 vss.n446 vss.n445 1245.36
R138 vss.n221 vss.n220 1058.82
R139 vss.n221 vss.n104 1058.82
R140 vss.n234 vss.n104 1058.82
R141 vss.n235 vss.n234 1058.82
R142 vss.n236 vss.n235 1058.82
R143 vss.n238 vss.n97 1058.82
R144 vss.n251 vss.n97 1058.82
R145 vss.n252 vss.n251 1058.82
R146 vss.n266 vss.n252 1058.82
R147 vss.n266 vss.n265 1058.82
R148 vss.n464 vss.t26 968.468
R149 vss.n265 vss.n264 951.085
R150 vss.n23 vss.n20 903.91
R151 vss.n449 vss.t26 783.348
R152 vss.n315 vss.n314 767.418
R153 vss.n236 vss.t0 717.648
R154 vss.t30 vss.n313 687.957
R155 vss.n307 vss.n306 635.574
R156 vss.n215 vss.n214 588.759
R157 vss.n218 vss.n111 588.759
R158 vss.n355 vss.n354 588.515
R159 vss.n255 vss.n96 585
R160 vss.n265 vss.n96 585
R161 vss.n268 vss.n267 585
R162 vss.n267 vss.n266 585
R163 vss.n95 vss.n93 585
R164 vss.n252 vss.n95 585
R165 vss.n250 vss.n249 585
R166 vss.n251 vss.n250 585
R167 vss.n99 vss.n98 585
R168 vss.n98 vss.n97 585
R169 vss.n240 vss.n239 585
R170 vss.n239 vss.n238 585
R171 vss.n237 vss.n102 585
R172 vss.n237 vss.n236 585
R173 vss.n107 vss.n103 585
R174 vss.n235 vss.n103 585
R175 vss.n233 vss.n232 585
R176 vss.n234 vss.n233 585
R177 vss.n224 vss.n105 585
R178 vss.n105 vss.n104 585
R179 vss.n223 vss.n222 585
R180 vss.n222 vss.n221 585
R181 vss.n219 vss.n109 585
R182 vss.n220 vss.n219 585
R183 vss.n213 vss.n117 585
R184 vss.n120 vss.n116 585
R185 vss.n217 vss.n116 585
R186 vss.n208 vss.n207 585
R187 vss.n200 vss.n123 585
R188 vss.n202 vss.n201 585
R189 vss.n193 vss.n125 585
R190 vss.n195 vss.n194 585
R191 vss.n186 vss.n182 585
R192 vss.n188 vss.n187 585
R193 vss.n184 vss.n110 585
R194 vss.n218 vss.n217 585
R195 vss.n254 vss.n253 585
R196 vss.n258 vss.n257 585
R197 vss.n83 vss.n81 585
R198 vss.n256 vss.n81 585
R199 vss.n276 vss.n275 585
R200 vss.n277 vss.n276 585
R201 vss.n87 vss.n79 585
R202 vss.n280 vss.n79 585
R203 vss.n282 vss.n80 585
R204 vss.n282 vss.n281 585
R205 vss.n287 vss.n286 585
R206 vss.n286 vss.n285 585
R207 vss.n78 vss.n76 585
R208 vss.n284 vss.n78 585
R209 vss.n72 vss.n69 585
R210 vss.n283 vss.n69 585
R211 vss.n295 vss.n294 585
R212 vss.n296 vss.n295 585
R213 vss.n70 vss.n68 585
R214 vss.n297 vss.n68 585
R215 vss.n299 vss.n60 585
R216 vss.n299 vss.n298 585
R217 vss.n263 vss.n262 585
R218 vss.n264 vss.n263 585
R219 vss.n301 vss.n300 585
R220 vss.n304 vss.n303 585
R221 vss.n143 vss.n62 585
R222 vss.n150 vss.n149 585
R223 vss.n148 vss.n142 585
R224 vss.n175 vss.n174 585
R225 vss.n173 vss.n172 585
R226 vss.n164 vss.n140 585
R227 vss.n166 vss.n165 585
R228 vss.n162 vss.n161 585
R229 vss.n160 vss.n159 585
R230 vss.n119 vss.n118 585
R231 vss.n448 vss.t47 576.794
R232 vss.n314 vss.t30 522.764
R233 vss.n355 vss.n353 512.625
R234 vss.t50 vss.t47 502.747
R235 vss.t51 vss.t50 502.747
R236 vss.t48 vss.t51 502.747
R237 vss.n431 vss.t65 493.086
R238 vss.n467 vss.t65 493.086
R239 vss.n264 vss.n253 435.913
R240 vss.n298 vss.n297 408.67
R241 vss.n297 vss.n296 408.67
R242 vss.n284 vss.n283 408.67
R243 vss.n285 vss.n284 408.67
R244 vss.n281 vss.n280 408.67
R245 vss.n257 vss.n256 408.67
R246 vss.n257 vss.n253 408.67
R247 vss.n431 vss.n430 391.663
R248 vss.n238 vss.t0 341.176
R249 vss.n442 vss.t0 314.589
R250 vss.n55 vss.t0 311.781
R251 vss.n436 vss.n426 307.036
R252 vss.n348 vss.n347 292.5
R253 vss.n347 vss.n346 292.5
R254 vss.n370 vss.n369 292.5
R255 vss.n369 vss.n368 292.5
R256 vss.n279 vss.t26 287.067
R257 vss.n308 vss.n30 281.336
R258 vss.n446 vss.n30 281.243
R259 vss.t1 vss.n441 279.022
R260 vss.n322 vss.n319 270.709
R261 vss.n256 vss.t0 267.906
R262 vss.n461 vss.n10 262.366
R263 vss.n226 vss.n108 258.334
R264 vss.n215 vss.n118 257.466
R265 vss.n436 vss.n435 256.805
R266 vss.n444 vss.n32 255.26
R267 vss.n217 vss.n216 254.34
R268 vss.n217 vss.n112 254.34
R269 vss.n217 vss.n113 254.34
R270 vss.n217 vss.n114 254.34
R271 vss.n217 vss.n115 254.34
R272 vss.n260 vss.n259 254.34
R273 vss.n306 vss.n59 254.34
R274 vss.n302 vss.n301 254.34
R275 vss.n301 vss.n67 254.34
R276 vss.n301 vss.n66 254.34
R277 vss.n301 vss.n65 254.34
R278 vss.n301 vss.n64 254.34
R279 vss.n301 vss.n63 254.34
R280 vss.n462 vss.n9 252.304
R281 vss.n296 vss.t0 249.743
R282 vss.n219 vss.n218 249.663
R283 vss.n368 vss.n318 232.525
R284 vss.n280 vss.n279 227.038
R285 vss.n451 vss.n27 223.468
R286 vss.n469 vss.n2 216.017
R287 vss.n281 vss.t0 213.417
R288 vss.n421 vss.n35 200.388
R289 vss.n442 vss.t28 199
R290 vss.n368 vss.n367 195.305
R291 vss.n285 vss.t0 195.254
R292 vss.n52 vss.n51 194.863
R293 vss.t25 vss.t24 191.542
R294 vss.n51 vss.t0 190.965
R295 vss.n400 vss.t36 189.031
R296 vss.n272 vss.n91 185
R297 vss.n274 vss.n273 185
R298 vss.n89 vss.n88 185
R299 vss.n86 vss.n85 185
R300 vss.n77 vss.n75 185
R301 vss.n289 vss.n288 185
R302 vss.n291 vss.n74 185
R303 vss.n293 vss.n292 185
R304 vss.n144 vss.n71 185
R305 vss.n145 vss.n61 185
R306 vss.n145 vss.t14 185
R307 vss.n147 vss.n146 185
R308 vss.n152 vss.n151 185
R309 vss.n153 vss.n139 185
R310 vss.n155 vss.n138 185
R311 vss.n171 vss.n170 185
R312 vss.n168 vss.n167 185
R313 vss.n163 vss.n156 185
R314 vss.n156 vss.t14 185
R315 vss.n158 vss.n157 185
R316 vss.n212 vss.n211 185
R317 vss.n210 vss.n209 185
R318 vss.n206 vss.n205 185
R319 vss.n204 vss.n203 185
R320 vss.n199 vss.n198 185
R321 vss.n197 vss.n196 185
R322 vss.n192 vss.n191 185
R323 vss.n190 vss.n189 185
R324 vss.n185 vss.n108 185
R325 vss.n270 vss.n269 185
R326 vss.n248 vss.n92 185
R327 vss.n247 vss.n246 185
R328 vss.n244 vss.n100 185
R329 vss.n242 vss.n241 185
R330 vss.n178 vss.n101 185
R331 vss.n231 vss.n230 185
R332 vss.n228 vss.n106 185
R333 vss.n226 vss.n225 185
R334 vss.n435 vss.n434 184.031
R335 vss.n279 vss.n277 181.631
R336 vss.n427 vss.n426 177.084
R337 vss.n117 vss.n116 175.546
R338 vss.n207 vss.n116 175.546
R339 vss.n201 vss.n200 175.546
R340 vss.n194 vss.n193 175.546
R341 vss.n187 vss.n186 175.546
R342 vss.n218 vss.n110 175.546
R343 vss.n161 vss.n160 175.546
R344 vss.n165 vss.n164 175.546
R345 vss.n174 vss.n173 175.546
R346 vss.n149 vss.n148 175.546
R347 vss.n303 vss.n62 175.546
R348 vss.n299 vss.n68 175.546
R349 vss.n295 vss.n68 175.546
R350 vss.n295 vss.n69 175.546
R351 vss.n78 vss.n69 175.546
R352 vss.n286 vss.n78 175.546
R353 vss.n286 vss.n282 175.546
R354 vss.n282 vss.n79 175.546
R355 vss.n276 vss.n79 175.546
R356 vss.n276 vss.n81 175.546
R357 vss.n258 vss.n81 175.546
R358 vss.n222 vss.n219 175.546
R359 vss.n222 vss.n105 175.546
R360 vss.n233 vss.n105 175.546
R361 vss.n233 vss.n103 175.546
R362 vss.n237 vss.n103 175.546
R363 vss.n239 vss.n237 175.546
R364 vss.n239 vss.n98 175.546
R365 vss.n250 vss.n98 175.546
R366 vss.n250 vss.n95 175.546
R367 vss.n267 vss.n95 175.546
R368 vss.n267 vss.n96 175.546
R369 vss.n263 vss.n96 175.546
R370 vss.n453 vss.n452 169.446
R371 vss.n145 vss.n144 163.333
R372 vss.n283 vss.t0 158.928
R373 vss.n302 vss.n59 152.643
R374 vss.n157 vss.n156 150
R375 vss.n168 vss.n156 150
R376 vss.n170 vss.n155 150
R377 vss.n153 vss.n152 150
R378 vss.n146 vss.n145 150
R379 vss.n211 vss.n210 150
R380 vss.n205 vss.n204 150
R381 vss.n198 vss.n197 150
R382 vss.n191 vss.n190 150
R383 vss.n230 vss.n228 150
R384 vss.n242 vss.n101 150
R385 vss.n246 vss.n244 150
R386 vss.n270 vss.n92 150
R387 vss.n292 vss.n291 150
R388 vss.n289 vss.n75 150
R389 vss.n89 vss.n85 150
R390 vss.n273 vss.n272 150
R391 vss.n348 vss.n342 149.538
R392 vss.n445 vss.n444 147.642
R393 vss.n300 vss.n299 146.287
R394 vss.t38 vss.n399 141.774
R395 vss.n277 vss.t0 140.764
R396 vss.n263 vss.n254 138.486
R397 vss.n420 vss.n36 137.462
R398 vss.n395 vss.n318 129.227
R399 vss.n342 vss.n332 126.4
R400 vss.n413 vss.n36 122.373
R401 vss.n404 vss.n46 113.549
R402 vss.t28 vss.t1 113.472
R403 vss.n441 vss.n440 111.778
R404 vss.n353 vss.n46 109.558
R405 vss.n373 vss.n331 104.918
R406 vss.n301 vss.t0 105.091
R407 vss.n298 vss.t0 104.439
R408 vss.n396 vss.t36 99.1166
R409 vss.n365 vss.n364 97.5005
R410 vss.n366 vss.n365 97.5005
R411 vss.n344 vss.n341 97.5005
R412 vss.n345 vss.n344 97.5005
R413 vss.n429 vss.n428 89.9525
R414 vss.n352 vss.t21 89.2211
R415 vss.n352 vss.t23 89.0687
R416 vss.t63 vss.t25 84.8974
R417 vss.t20 vss.n343 84.4265
R418 vss.n343 vss.t22 82.5503
R419 vss.n310 vss.n309 76.8967
R420 vss.n345 vss.t20 76.4529
R421 vss.n216 vss.n215 76.3222
R422 vss.n207 vss.n112 76.3222
R423 vss.n201 vss.n113 76.3222
R424 vss.n194 vss.n114 76.3222
R425 vss.n187 vss.n115 76.3222
R426 vss.n160 vss.n63 76.3222
R427 vss.n165 vss.n64 76.3222
R428 vss.n173 vss.n65 76.3222
R429 vss.n148 vss.n66 76.3222
R430 vss.n67 vss.n62 76.3222
R431 vss.n300 vss.n59 76.3222
R432 vss.n259 vss.n254 76.3222
R433 vss.n216 vss.n117 76.3222
R434 vss.n200 vss.n112 76.3222
R435 vss.n193 vss.n113 76.3222
R436 vss.n186 vss.n114 76.3222
R437 vss.n115 vss.n110 76.3222
R438 vss.n259 vss.n258 76.3222
R439 vss.n303 vss.n302 76.3222
R440 vss.n149 vss.n67 76.3222
R441 vss.n174 vss.n66 76.3222
R442 vss.n164 vss.n65 76.3222
R443 vss.n161 vss.n64 76.3222
R444 vss.n118 vss.n63 76.3222
R445 vss.n211 vss.n121 74.5978
R446 vss.n157 vss.n121 74.5978
R447 vss.n56 vss.n55 74.0483
R448 vss.n341 vss.n340 73.0981
R449 vss.n271 vss.n270 69.3109
R450 vss.n272 vss.n271 69.3109
R451 vss.n27 vss.n9 69.0601
R452 vss.n90 vss.t14 65.8183
R453 vss.n84 vss.t14 65.8183
R454 vss.n290 vss.t14 65.8183
R455 vss.t14 vss.n73 65.8183
R456 vss.n141 vss.t14 65.8183
R457 vss.n154 vss.t14 65.8183
R458 vss.n169 vss.t14 65.8183
R459 vss.n122 vss.t14 65.8183
R460 vss.n124 vss.t14 65.8183
R461 vss.n126 vss.t14 65.8183
R462 vss.n183 vss.t14 65.8183
R463 vss.n245 vss.t14 65.8183
R464 vss.n243 vss.t14 65.8183
R465 vss.n229 vss.t14 65.8183
R466 vss.n227 vss.t14 65.8183
R467 vss.n313 vss.t26 65.4995
R468 vss.n350 vss.n339 65.0005
R469 vss.n343 vss.n339 65.0005
R470 vss.n340 vss.n338 65.0005
R471 vss.n343 vss.n338 65.0005
R472 vss.n309 vss.n308 65.0005
R473 vss.n447 vss.n446 65.0005
R474 vss.n448 vss.n447 65.0005
R475 vss.t0 vss.t48 60.4079
R476 vss.t10 vss.t0 60.4079
R477 vss.t53 vss.t0 60.4079
R478 vss.n271 vss.t14 57.8461
R479 vss.n52 vss.t10 56.5107
R480 vss.n56 vss.t53 56.5107
R481 vss.n364 vss.n340 56.241
R482 vss.n121 vss.t14 55.2026
R483 vss.n18 vss.n13 54.0035
R484 vss.n16 vss.n14 54.0035
R485 vss.n407 vss.n43 53.9338
R486 vss.n409 vss.n42 53.9338
R487 vss.n169 vss.n168 53.3664
R488 vss.n155 vss.n154 53.3664
R489 vss.n152 vss.n141 53.3664
R490 vss.n210 vss.n122 53.3664
R491 vss.n204 vss.n124 53.3664
R492 vss.n197 vss.n126 53.3664
R493 vss.n190 vss.n183 53.3664
R494 vss.n227 vss.n226 53.3664
R495 vss.n230 vss.n229 53.3664
R496 vss.n243 vss.n242 53.3664
R497 vss.n246 vss.n245 53.3664
R498 vss.n292 vss.n73 53.3664
R499 vss.n290 vss.n289 53.3664
R500 vss.n85 vss.n84 53.3664
R501 vss.n273 vss.n90 53.3664
R502 vss.n90 vss.n89 53.3664
R503 vss.n84 vss.n75 53.3664
R504 vss.n291 vss.n290 53.3664
R505 vss.n144 vss.n73 53.3664
R506 vss.n146 vss.n141 53.3664
R507 vss.n154 vss.n153 53.3664
R508 vss.n170 vss.n169 53.3664
R509 vss.n205 vss.n122 53.3664
R510 vss.n198 vss.n124 53.3664
R511 vss.n191 vss.n126 53.3664
R512 vss.n183 vss.n108 53.3664
R513 vss.n245 vss.n92 53.3664
R514 vss.n244 vss.n243 53.3664
R515 vss.n229 vss.n101 53.3664
R516 vss.n228 vss.n227 53.3664
R517 vss.n4 vss.n1 53.1823
R518 vss.t65 vss.n4 53.1823
R519 vss.n3 vss.n2 53.1823
R520 vss.t65 vss.n3 53.1823
R521 vss.t0 vss.t49 53.1497
R522 vss.t0 vss.t15 53.1497
R523 vss.t0 vss.t19 53.1497
R524 vss.t0 vss.t16 53.1497
R525 vss.t0 vss.t17 53.1497
R526 vss.t0 vss.t11 53.1497
R527 vss.t0 vss.t9 53.1497
R528 vss.t0 vss.t12 53.1497
R529 vss.t0 vss.t13 53.1497
R530 vss.t0 vss.t54 53.1497
R531 vss.t0 vss.t56 53.1497
R532 vss.t0 vss.t52 53.1497
R533 vss.t0 vss.t55 53.1497
R534 vss.n399 vss.n315 49.7676
R535 vss.n402 vss.n401 48.7505
R536 vss.n401 vss.n400 48.7505
R537 vss.n394 vss.n393 48.7505
R538 vss.n395 vss.n394 48.7505
R539 vss.n366 vss.t5 45.4967
R540 vss.n311 vss.n310 44.185
R541 vss.n470 vss.n469 42.0571
R542 vss.n435 vss.n2 41.1681
R543 vss.n367 vss.n366 39.8683
R544 vss.n22 vss.n21 39.7638
R545 vss.n453 vss.n24 39.511
R546 vss.n278 vss.t18 39.3863
R547 vss.n342 vss.n335 34.4123
R548 vss.t5 vss.n335 34.4123
R549 vss.n351 vss.n334 34.4123
R550 vss.t5 vss.n334 34.4123
R551 vss.n469 vss.n468 34.4123
R552 vss.n468 vss.n467 34.4123
R553 vss.n433 vss.n432 34.4123
R554 vss.n432 vss.n431 34.4123
R555 vss.n404 vss.n403 33.9329
R556 vss.n326 vss.n50 32.5005
R557 vss.t63 vss.n50 32.5005
R558 vss.n375 vss.n49 32.5005
R559 vss.t63 vss.n49 32.5005
R560 vss.n22 vss.n8 32.5005
R561 vss.n440 vss.n8 32.5005
R562 vss.n27 vss.n7 32.5005
R563 vss.n314 vss.n7 32.5005
R564 vss.t22 vss.t5 32.3638
R565 vss.n421 vss.n420 32.1396
R566 vss.n1 vss.t66 30.8834
R567 vss.n363 vss.n333 30.4707
R568 vss.n346 vss.n345 28.6115
R569 vss.n326 vss.n320 28.0594
R570 vss.n130 vss.t7 26.6016
R571 vss.n37 vss.t39 25.1357
R572 vss.n376 vss.n374 24.7516
R573 vss.n403 vss.n47 24.4644
R574 vss.n445 vss.n31 23.8095
R575 vss.n308 vss.n307 23.4151
R576 vss.n428 vss.n427 23.0405
R577 vss.n135 vss.n127 20.7857
R578 vss.n134 vss.n128 20.7857
R579 vss.n130 vss.n129 20.7857
R580 vss.n411 vss.n41 20.7665
R581 vss.n412 vss.n40 20.7665
R582 vss.n415 vss.n39 20.7665
R583 vss.n416 vss.n38 20.7665
R584 vss.n349 vss.n348 20.517
R585 vss.n397 vss.n47 20.1729
R586 vss.n397 vss.n396 20.1729
R587 vss.n356 vss.n316 20.1729
R588 vss.n396 vss.n316 20.1729
R589 vss.n349 vss.n341 20.0772
R590 vss.n388 vss.n387 19.4026
R591 vss.t24 vss.n395 19.2382
R592 vss.n392 vss.n320 19.2005
R593 vss.n398 vss.n46 18.8715
R594 vss.n399 vss.n398 18.8715
R595 vss.n354 vss.n317 18.8715
R596 vss.n318 vss.n317 18.8715
R597 vss.n433 vss.n429 18.7337
R598 vss.n307 vss.n58 17.5097
R599 vss.n374 vss.n319 17.1218
R600 vss.n387 vss.n48 16.4046
R601 vss.n434 vss.n433 16.3845
R602 vss.n403 vss.n402 16.1396
R603 vss.n132 vss.n131 16.0068
R604 vss.n462 vss.n461 15.5385
R605 vss.n422 vss.n421 14.6255
R606 vss.n442 vss.n422 14.6255
R607 vss.n444 vss.n443 14.6255
R608 vss.n443 vss.n442 14.6255
R609 vss.n329 vss.n328 14.0913
R610 vss.n387 vss.n386 12.7191
R611 vss.n279 vss.n278 12.1537
R612 vss.n434 vss.n425 11.9393
R613 vss.n430 vss.n425 11.9393
R614 vss.n426 vss.n424 11.9393
R615 vss.n424 vss.n5 11.9393
R616 vss.n43 vss.t35 11.6005
R617 vss.n43 vss.t32 11.6005
R618 vss.n42 vss.t27 11.6005
R619 vss.n42 vss.t29 11.6005
R620 vss.n13 vss.t33 11.6005
R621 vss.n13 vss.t34 11.6005
R622 vss.n14 vss.t31 11.6005
R623 vss.n14 vss.t37 11.6005
R624 vss.n452 vss.n451 10.5495
R625 vss.n429 vss.n1 10.0532
R626 vss.n371 vss.n333 9.74099
R627 vss.n390 vss.n322 9.3005
R628 vss.n454 vss.n453 9.3005
R629 vss.n459 vss.n10 9.3005
R630 vss.n20 vss.n12 9.3005
R631 vss.n350 vss.n349 8.86924
R632 vss.n370 vss.n332 8.42977
R633 vss.n396 vss.t63 7.5283
R634 vss.n427 vss.n423 7.5005
R635 vss.n438 vss.n423 7.5005
R636 vss.n437 vss.n436 7.5005
R637 vss.n438 vss.n437 7.5005
R638 vss.n376 vss.n375 7.34725
R639 vss.n373 vss.n372 7.32557
R640 vss.n31 vss.n29 7.313
R641 vss.n51 vss.n29 7.313
R642 vss.n30 vss.n28 7.313
R643 vss.n51 vss.n28 7.313
R644 vss.n374 vss.n373 6.9983
R645 vss.n420 vss.n419 6.9005
R646 vss.n418 vss.n36 6.9005
R647 vss.n385 vss 6.21282
R648 vss.n58 vss.n33 6.15839
R649 vss.n55 vss.n33 6.15839
R650 vss.n34 vss.n32 6.15839
R651 vss.n441 vss.n34 6.15839
R652 vss.n363 vss.n362 5.92892
R653 vss.n372 vss.n371 5.77749
R654 vss.n351 vss.n350 5.73359
R655 vss.n364 vss.n363 5.34506
R656 vss.n278 vss.t0 4.95804
R657 vss.n159 vss.n119 4.90263
R658 vss.n223 vss.n109 4.90263
R659 vss.n451 vss.n450 4.8755
R660 vss.n450 vss.n449 4.8755
R661 vss.n463 vss.n462 4.8755
R662 vss.n464 vss.n463 4.8755
R663 vss.n225 vss.n223 4.84816
R664 vss.n224 vss.n106 4.84816
R665 vss.n232 vss.n231 4.84816
R666 vss.n241 vss.n102 4.84816
R667 vss.n240 vss.n100 4.84816
R668 vss.n247 vss.n99 4.84816
R669 vss.n249 vss.n248 4.84816
R670 vss.n269 vss.n93 4.84816
R671 vss.n262 vss.n255 4.57193
R672 vss.n454 vss.n26 4.5005
R673 vss.n386 vss.n385 4.5005
R674 vss.n45 vss.n44 4.5005
R675 vss.n390 vss.n323 4.5005
R676 vss.n459 vss.n458 4.5005
R677 vss.n457 vss.n12 4.5005
R678 vss.n41 vss.t4 4.3505
R679 vss.n41 vss.t43 4.3505
R680 vss.n40 vss.t2 4.3505
R681 vss.n40 vss.t46 4.3505
R682 vss.n39 vss.t3 4.3505
R683 vss.n39 vss.t8 4.3505
R684 vss.n38 vss.t57 4.3505
R685 vss.n38 vss.t62 4.3505
R686 vss.n127 vss.t42 4.3505
R687 vss.n127 vss.t44 4.3505
R688 vss.n128 vss.t45 4.3505
R689 vss.n128 vss.t60 4.3505
R690 vss.n129 vss.t40 4.3505
R691 vss.n129 vss.t59 4.3505
R692 vss.n457 vss.n0 4.26937
R693 vss.n15 vss.n11 4.25229
R694 vss.n460 vss.n459 4.1668
R695 vss.n419 vss.n37 4.10351
R696 vss.n16 vss.n15 4.02718
R697 vss.n407 vss.n406 3.98965
R698 vss.n354 vss.n331 3.98739
R699 vss.n260 vss.n35 3.9624
R700 vss.n159 vss.n158 3.81327
R701 vss.n163 vss.n162 3.81327
R702 vss.n167 vss.n166 3.81327
R703 vss.n171 vss.n140 3.81327
R704 vss.n172 vss.n138 3.81327
R705 vss.n175 vss.n139 3.81327
R706 vss.n151 vss.n142 3.81327
R707 vss.n150 vss.n147 3.81327
R708 vss.n143 vss.n61 3.81327
R709 vss.n21 vss.n10 3.76521
R710 vss.n470 vss.n1 3.71562
R711 vss.n255 vss.n94 3.55606
R712 vss.n179 vss.n178 3.48646
R713 vss.n471 vss.n0 3.33015
R714 vss.n328 vss.t67 3.16414
R715 vss.n328 vss.t64 3.16414
R716 vss.n15 vss.n9 3.10035
R717 vss.n388 vss.n326 2.96471
R718 vss.n217 vss.t0 128.062
R719 vss.n213 vss.n212 2.7239
R720 vss.n209 vss.n120 2.7239
R721 vss.n208 vss.n206 2.7239
R722 vss.n203 vss.n123 2.7239
R723 vss.n202 vss.n199 2.7239
R724 vss.n195 vss.n192 2.7239
R725 vss.n189 vss.n182 2.7239
R726 vss.n188 vss.n185 2.7239
R727 vss.n358 vss.n357 2.68591
R728 vss.n400 vss.t38 2.50977
R729 vss.n360 vss.n333 2.3255
R730 vss.n454 vss.n25 2.29617
R731 vss.n419 vss.n418 2.28754
R732 vss.n456 vss.n19 2.24795
R733 vss.n212 vss.n120 2.17922
R734 vss.n209 vss.n208 2.17922
R735 vss.n206 vss.n123 2.17922
R736 vss.n203 vss.n202 2.17922
R737 vss.n199 vss.n125 2.17922
R738 vss.n196 vss.n195 2.17922
R739 vss.n192 vss.n182 2.17922
R740 vss.n189 vss.n188 2.17922
R741 vss.n185 vss.n184 2.17922
R742 vss.n70 vss.n60 2.17819
R743 vss.n17 vss.n16 2.15904
R744 vss.n458 vss.n18 2.12067
R745 vss.n357 vss.n353 2.10102
R746 vss.n136 vss.n82 1.89157
R747 vss.n294 vss.n71 1.79105
R748 vss.n293 vss.n72 1.79105
R749 vss.n76 vss.n74 1.79105
R750 vss.n288 vss.n287 1.79105
R751 vss.n80 vss.n77 1.79105
R752 vss.n274 vss.n83 1.79105
R753 vss.n18 vss.n17 1.78099
R754 vss.n471 vss.n470 1.7255
R755 vss.n131 vss 1.7155
R756 vss.n181 vss.n125 1.68901
R757 vss.n411 vss.n410 1.67152
R758 vss.n306 vss.n305 1.64587
R759 vss.n312 vss.t0 1.63432
R760 vss.n359 vss.n358 1.55732
R761 vss.n180 vss.n179 1.51978
R762 vss.n362 vss.n351 1.47378
R763 vss.n135 vss.n134 1.46641
R764 vss.n133 vss.n130 1.43989
R765 vss.n87 vss 1.37971
R766 vss.n91 vss.n35 1.37971
R767 vss.n310 vss.t0 1.37561
R768 vss.n179 vss.n107 1.3622
R769 vss.n24 vss.n23 1.30961
R770 vss.n408 vss.n407 1.23783
R771 vss.n275 vss.n82 1.18613
R772 vss.n410 vss.n409 1.13184
R773 vss.n261 vss.n260 1.11796
R774 vss.n162 vss.n158 1.08986
R775 vss.n166 vss.n163 1.08986
R776 vss.n167 vss.n140 1.08986
R777 vss.n172 vss.n171 1.08986
R778 vss.n142 vss.n139 1.08986
R779 vss.n151 vss.n150 1.08986
R780 vss.n147 vss.n143 1.08986
R781 vss.n304 vss.n61 1.08986
R782 vss.n305 vss.n304 1.08986
R783 vss.n268 vss.n94 1.08986
R784 vss.t61 vss.t41 1.07946
R785 vss.n439 vss.n438 1.07946
R786 vss.t58 vss.t6 1.07946
R787 vss.n406 vss.n44 1.07186
R788 vss.n23 vss.n22 1.06085
R789 vss.n405 vss.n45 1.05279
R790 vss.n196 vss.n181 1.03539
R791 vss.n405 vss.n404 1.03383
R792 vss.n412 vss.n411 0.998567
R793 vss.n416 vss.n415 0.997923
R794 vss.n409 vss.n408 0.995892
R795 vss.n176 vss.n138 0.871989
R796 vss.n214 vss.n119 0.817521
R797 vss.n111 vss.n109 0.817521
R798 vss.n305 vss.n60 0.798988
R799 vss.n322 vss.n320 0.775237
R800 vss.n180 vss.n177 0.765632
R801 vss.n132 vss.n58 0.739443
R802 vss.n21 vss.n20 0.684992
R803 vss.n375 vss.n47 0.682157
R804 vss.n177 vss.n137 0.653909
R805 vss.n417 vss.n416 0.633876
R806 vss.n88 vss.n82 0.605415
R807 vss.n181 vss.n180 0.596304
R808 vss.n177 vss.n176 0.59175
R809 vss.n137 vss.n135 0.539326
R810 vss.n413 vss.n32 0.532356
R811 vss.n414 vss.n412 0.528206
R812 vss.n390 vss.n389 0.47062
R813 vss.n415 vss.n414 0.469572
R814 vss.n455 vss.n454 0.469344
R815 vss.n324 vss.n323 0.456098
R816 vss.n137 vss.n136 0.452967
R817 vss.n379 vss.n377 0.452003
R818 vss.n406 vss.n405 0.4505
R819 vss.n455 vss.n12 0.441368
R820 vss vss.n86 0.411842
R821 vss.n323 vss.n321 0.399345
R822 vss.n357 vss.n356 0.391918
R823 vss.n71 vss.n70 0.387646
R824 vss.n294 vss.n293 0.387646
R825 vss.n74 vss.n72 0.387646
R826 vss.n288 vss.n76 0.387646
R827 vss.n287 vss.n77 0.387646
R828 vss.n88 vss.n87 0.387646
R829 vss.n275 vss.n274 0.387646
R830 vss.n91 vss.n83 0.387646
R831 vss.n377 vss.n330 0.376108
R832 vss.n360 vss.n359 0.368932
R833 vss.n361 vss.n360 0.355
R834 vss.n389 vss.n325 0.350102
R835 vss.n327 vss.n324 0.344129
R836 vss.n418 vss.n417 0.343093
R837 vss.n455 vss.n24 0.32741
R838 vss.n214 vss.n213 0.327309
R839 vss.n379 vss.n378 0.326722
R840 vss.n457 vss.n456 0.317677
R841 vss.n330 vss.n321 0.312188
R842 vss.n358 vss.n331 0.3005
R843 vss.n391 vss.n390 0.272145
R844 vss vss.n80 0.242466
R845 vss.n384 vss.n383 0.226831
R846 vss.n393 vss.n319 0.224276
R847 vss.n392 vss.n391 0.221929
R848 vss.n380 vss.n379 0.221128
R849 vss.n382 vss.n325 0.220839
R850 vss.n176 vss.n175 0.218372
R851 vss.n378 vss.n329 0.216846
R852 vss.n381 vss.n380 0.20954
R853 vss.n131 vss.n31 0.188367
R854 vss.n371 vss.n370 0.187817
R855 vss.n356 vss.n355 0.180782
R856 vss.n86 vss 0.14568
R857 vss.n428 vss.n0 0.139042
R858 vss.n381 vss.n48 0.133357
R859 vss.n377 vss.n376 0.126176
R860 vss.n456 vss.n455 0.1255
R861 vss.n362 vss.n361 0.122868
R862 vss vss.n471 0.120187
R863 vss.n361 vss.n352 0.118284
R864 vss.n184 vss.n111 0.109436
R865 vss.n389 vss.n388 0.107397
R866 vss.n133 vss.n132 0.0987955
R867 vss.n136 vss.n37 0.0948141
R868 vss.n19 vss 0.0874816
R869 vss.n410 vss.n26 0.0851774
R870 vss.n461 vss.n460 0.0850455
R871 vss.n417 vss 0.0849072
R872 vss.n414 vss.n413 0.0736577
R873 vss.n459 vss.n12 0.0711522
R874 vss.n383 vss.n382 0.0605
R875 vss.n225 vss.n224 0.0549681
R876 vss.n232 vss.n106 0.0549681
R877 vss.n231 vss.n107 0.0549681
R878 vss.n178 vss.n102 0.0549681
R879 vss.n241 vss.n240 0.0549681
R880 vss.n100 vss.n99 0.0549681
R881 vss.n249 vss.n247 0.0549681
R882 vss.n248 vss.n93 0.0549681
R883 vss.n269 vss.n268 0.0549681
R884 vss.n262 vss.n261 0.0512937
R885 vss vss.n384 0.048119
R886 vss.n389 vss.n324 0.0459545
R887 vss.n393 vss.n392 0.0452552
R888 vss.n385 vss.n327 0.0448787
R889 vss.n386 vss.n325 0.0428729
R890 vss.n359 vss.n330 0.0382747
R891 vss.n17 vss.n11 0.0367903
R892 vss.n378 vss.n44 0.0330444
R893 vss.n380 vss.n45 0.0294548
R894 vss.n452 vss.n25 0.0286818
R895 vss.n134 vss.n133 0.0270152
R896 vss.n402 vss.n48 0.027001
R897 vss.n458 vss.n457 0.0246098
R898 vss.n26 vss.n19 0.0195092
R899 vss.n460 vss.n11 0.0135435
R900 vss.n408 vss.n25 0.0126951
R901 vss.n391 vss.n321 0.00969913
R902 vss.n384 vss.n327 0.00493787
R903 vss.n383 vss.n329 0.00234911
R904 vss.n382 vss.n381 0.00191243
R905 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 935.75
R906 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 235.982
R907 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 235.978
R908 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 190.305
R909 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 190.305
R910 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 190.305
R911 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 190.305
R912 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 190.305
R913 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 190.305
R914 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 95.3928
R915 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 95.3648
R916 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 95.1789
R917 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 95.1648
R918 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 95.1542
R919 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 95.1535
R920 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 94.8314
R921 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 94.8314
R922 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 94.8314
R923 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 94.8314
R924 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 94.8314
R925 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 94.8314
R926 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 94.8314
R927 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 94.8314
R928 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 94.8314
R929 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 94.8314
R930 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 94.8314
R931 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 94.8314
R932 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 94.8314
R933 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 94.8314
R934 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 94.8314
R935 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 94.8314
R936 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 94.8314
R937 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 94.8314
R938 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 94.8314
R939 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 94.8314
R940 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 94.8314
R941 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 94.8314
R942 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 94.8314
R943 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 84.0884
R944 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 83.5719
R945 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 83.5719
R946 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 83.5719
R947 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 83.5719
R948 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 73.19
R949 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 26.074
R950 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 26.074
R951 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 26.074
R952 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 25.7843
R953 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 10.2822
R954 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 9.66398
R955 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R956 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R957 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R958 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R959 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 9.3005
R960 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 9.3005
R961 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R962 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R963 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 9.3005
R964 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R965 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R966 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R967 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 9.3005
R968 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R969 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R970 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R971 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 9.3005
R972 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R973 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R974 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R975 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R976 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 9.3005
R977 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 9.3005
R978 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 9.3005
R979 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 9.3005
R980 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 9.3005
R981 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 9.3005
R982 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 9.3005
R983 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 7.22993
R984 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 7.22993
R985 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 7.22993
R986 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 6.83022
R987 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 6.81633
R988 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 6.81633
R989 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 6.81633
R990 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 6.75312
R991 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 4.64588
R992 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 4.64588
R993 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 4.64588
R994 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 4.64588
R995 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 2.29815
R996 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 1.86108
R997 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 1.86108
R998 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 1.86108
R999 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 1.86108
R1000 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 1.86108
R1001 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 1.86108
R1002 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 1.86108
R1003 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 1.28692
R1004 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 1.25468
R1005 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 1.14402
R1006 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 1.1424
R1007 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 1.12066
R1008 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 1.12066
R1009 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 1.11251
R1010 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 1.10979
R1011 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 1.10164
R1012 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 1.10164
R1013 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 1.10164
R1014 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 1.10164
R1015 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 1.09892
R1016 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 1.09349
R1017 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 1.09349
R1018 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 1.08805
R1019 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 1.08262
R1020 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 1.08262
R1021 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 1.08262
R1022 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 1.07024
R1023 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 1.0237
R1024 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.959578
R1025 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 0.812055
R1026 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.77514
R1027 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.701365
R1028 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.645119
R1029 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 0.645119
R1030 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 0.645119
R1031 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 0.645119
R1032 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 0.645119
R1033 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 0.645119
R1034 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 0.645119
R1035 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.645119
R1036 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 0.645119
R1037 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.645119
R1038 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 0.645119
R1039 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 0.645119
R1040 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 0.645119
R1041 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 0.645119
R1042 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 0.645119
R1043 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.645119
R1044 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 0.645119
R1045 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.645119
R1046 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 0.645119
R1047 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 0.645119
R1048 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 0.645119
R1049 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 0.645119
R1050 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 0.645119
R1051 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.645119
R1052 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.645119
R1053 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 0.645119
R1054 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 0.645119
R1055 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 0.645119
R1056 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 0.645119
R1057 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 0.645118
R1058 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 0.590702
R1059 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 0.572258
R1060 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 0.495065
R1061 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.495065
R1062 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 0.481478
R1063 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.481478
R1064 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.475521
R1065 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 0.470609
R1066 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.470609
R1067 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 0.465174
R1068 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 0.465174
R1069 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.465174
R1070 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.459844
R1071 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 0.459739
R1072 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.459739
R1073 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 0.446152
R1074 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.446152
R1075 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.445943
R1076 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.443435
R1077 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.440717
R1078 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 0.440717
R1079 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.434551
R1080 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 0.432263
R1081 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.414484
R1082 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.408265
R1083 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.408265
R1084 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.40372
R1085 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.40372
R1086 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.314045
R1087 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 0.290206
R1088 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.0183279
R1089 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 0.0112346
R1090 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 0.0112346
R1091 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 0.0112346
R1092 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 0.0112346
R1093 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n93 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 0.0112346
R1094 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 0.0112346
R1095 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 0.0112346
R1096 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 0.0112346
R1097 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 0.00759293
R1098 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 0.00316393
R1099 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.t32 88.7532
R1100 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 22.2005
R1101 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 21.8665
R1102 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 21.5445
R1103 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 21.5445
R1104 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 21.5445
R1105 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 21.5445
R1106 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 21.5445
R1107 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 21.5445
R1108 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 21.5445
R1109 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 21.5445
R1110 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 21.5445
R1111 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 21.5445
R1112 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 21.5445
R1113 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 21.5445
R1114 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 21.5445
R1115 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 21.5418
R1116 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 4.3505
R1117 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 4.3505
R1118 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 4.3505
R1119 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 4.3505
R1120 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 4.3505
R1121 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 4.3505
R1122 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 4.3505
R1123 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 4.3505
R1124 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 4.3505
R1125 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 4.3505
R1126 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 4.3505
R1127 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 4.3505
R1128 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 4.3505
R1129 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 4.3505
R1130 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 4.3505
R1131 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 4.3505
R1132 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 4.3505
R1133 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 4.3505
R1134 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 4.3505
R1135 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 4.3505
R1136 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 4.3505
R1137 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 4.3505
R1138 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 4.3505
R1139 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 4.3505
R1140 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 4.3505
R1141 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 4.3505
R1142 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 4.3505
R1143 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 4.3505
R1144 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 4.3505
R1145 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 4.3505
R1146 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 4.3505
R1147 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 OTA_vref_0.OTA_vref_stage2_0.vref0.t0 4.3505
R1148 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 4.27517
R1149 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 3.08331
R1150 a_n1236_n9479.n58 a_n1236_n9479.t8 190.305
R1151 a_n1236_n9479.t8 a_n1236_n9479.n57 190.305
R1152 a_n1236_n9479.t26 a_n1236_n9479.n42 190.305
R1153 a_n1236_n9479.n56 a_n1236_n9479.t26 190.305
R1154 a_n1236_n9479.n23 a_n1236_n9479.t16 190.305
R1155 a_n1236_n9479.n21 a_n1236_n9479.t16 190.305
R1156 a_n1236_n9479.t30 a_n1236_n9479.n18 190.305
R1157 a_n1236_n9479.n20 a_n1236_n9479.t30 190.305
R1158 a_n1236_n9479.t12 a_n1236_n9479.n77 190.305
R1159 a_n1236_n9479.n81 a_n1236_n9479.t12 190.305
R1160 a_n1236_n9479.t22 a_n1236_n9479.n79 190.305
R1161 a_n1236_n9479.n80 a_n1236_n9479.t22 190.305
R1162 a_n1236_n9479.t10 a_n1236_n9479.n47 190.305
R1163 a_n1236_n9479.n48 a_n1236_n9479.t10 190.305
R1164 a_n1236_n9479.t24 a_n1236_n9479.n45 190.305
R1165 a_n1236_n9479.n49 a_n1236_n9479.t24 190.305
R1166 a_n1236_n9479.t28 a_n1236_n9479.n28 190.305
R1167 a_n1236_n9479.n32 a_n1236_n9479.t28 190.305
R1168 a_n1236_n9479.t2 a_n1236_n9479.n30 190.305
R1169 a_n1236_n9479.n31 a_n1236_n9479.t2 190.305
R1170 a_n1236_n9479.t18 a_n1236_n9479.n70 190.305
R1171 a_n1236_n9479.n71 a_n1236_n9479.t18 190.305
R1172 a_n1236_n9479.n16 a_n1236_n9479.t6 190.305
R1173 a_n1236_n9479.t6 a_n1236_n9479.n13 190.305
R1174 a_n1236_n9479.t20 a_n1236_n9479.n62 190.305
R1175 a_n1236_n9479.n63 a_n1236_n9479.t20 190.305
R1176 a_n1236_n9479.t4 a_n1236_n9479.n37 190.305
R1177 a_n1236_n9479.n64 a_n1236_n9479.t4 190.305
R1178 a_n1236_n9479.n25 a_n1236_n9479.t14 95.1811
R1179 a_n1236_n9479.n41 a_n1236_n9479.t0 95.1783
R1180 a_n1236_n9479.n54 a_n1236_n9479.n53 22.3176
R1181 a_n1236_n9479.n36 a_n1236_n9479.n35 22.2301
R1182 a_n1236_n9479.n9 a_n1236_n9479.n26 22.2284
R1183 a_n1236_n9479.n0 a_n1236_n9479.n27 22.2284
R1184 a_n1236_n9479.n6 a_n1236_n9479.n34 22.2284
R1185 a_n1236_n9479.n12 a_n1236_n9479.n69 22.2284
R1186 a_n1236_n9479.n68 a_n1236_n9479.n67 22.2284
R1187 a_n1236_n9479.n10 a_n1236_n9479.n38 22.2284
R1188 a_n1236_n9479.n40 a_n1236_n9479.n39 22.2284
R1189 a_n1236_n9479.n5 a_n1236_n9479.n17 22.1884
R1190 a_n1236_n9479.n1 a_n1236_n9479.n83 22.1884
R1191 a_n1236_n9479.n3 a_n1236_n9479.n43 22.1884
R1192 a_n1236_n9479.n2 a_n1236_n9479.n44 22.1884
R1193 a_n1236_n9479.n11 a_n1236_n9479.n51 22.1884
R1194 a_n1236_n9479.n8 a_n1236_n9479.n52 22.1884
R1195 a_n1236_n9479.n84 a_n1236_n9479.n4 22.1884
R1196 a_n1236_n9479.n59 a_n1236_n9479.n41 11.5566
R1197 a_n1236_n9479.n25 a_n1236_n9479.n24 10.9335
R1198 a_n1236_n9479.n77 a_n1236_n9479.n76 9.89233
R1199 a_n1236_n9479.n47 a_n1236_n9479.n15 9.89233
R1200 a_n1236_n9479.n24 a_n1236_n9479.n23 9.80925
R1201 a_n1236_n9479.n59 a_n1236_n9479.n58 9.80925
R1202 a_n1236_n9479.n64 a_n1236_n9479.n60 9.48127
R1203 a_n1236_n9479.n75 a_n1236_n9479.n13 9.40378
R1204 a_n1236_n9479.n31 a_n1236_n9479.n14 9.39819
R1205 a_n1236_n9479.n41 a_n1236_n9479.n40 4.9275
R1206 a_n1236_n9479.n9 a_n1236_n9479.n25 4.79654
R1207 a_n1236_n9479.n61 a_n1236_n9479.n10 4.5005
R1208 a_n1236_n9479.n66 a_n1236_n9479.n65 4.5005
R1209 a_n1236_n9479.n12 a_n1236_n9479.n72 4.5005
R1210 a_n1236_n9479.n74 a_n1236_n9479.n73 4.5005
R1211 a_n1236_n9479.n6 a_n1236_n9479.n33 4.5005
R1212 a_n1236_n9479.n29 a_n1236_n9479.n0 4.5005
R1213 a_n1236_n9479.n8 a_n1236_n9479.n7 4.5005
R1214 a_n1236_n9479.n55 a_n1236_n9479.n54 4.5005
R1215 a_n1236_n9479.n11 a_n1236_n9479.n50 4.5005
R1216 a_n1236_n9479.n46 a_n1236_n9479.n2 4.5005
R1217 a_n1236_n9479.n78 a_n1236_n9479.n3 4.5005
R1218 a_n1236_n9479.n1 a_n1236_n9479.n82 4.5005
R1219 a_n1236_n9479.n22 a_n1236_n9479.n5 4.5005
R1220 a_n1236_n9479.n19 a_n1236_n9479.n4 4.5005
R1221 a_n1236_n9479.n17 a_n1236_n9479.t37 4.3505
R1222 a_n1236_n9479.n17 a_n1236_n9479.t17 4.3505
R1223 a_n1236_n9479.n83 a_n1236_n9479.t35 4.3505
R1224 a_n1236_n9479.n83 a_n1236_n9479.t13 4.3505
R1225 a_n1236_n9479.n43 a_n1236_n9479.t23 4.3505
R1226 a_n1236_n9479.n43 a_n1236_n9479.t47 4.3505
R1227 a_n1236_n9479.n44 a_n1236_n9479.t34 4.3505
R1228 a_n1236_n9479.n44 a_n1236_n9479.t11 4.3505
R1229 a_n1236_n9479.n51 a_n1236_n9479.t25 4.3505
R1230 a_n1236_n9479.n51 a_n1236_n9479.t32 4.3505
R1231 a_n1236_n9479.n52 a_n1236_n9479.t43 4.3505
R1232 a_n1236_n9479.n52 a_n1236_n9479.t9 4.3505
R1233 a_n1236_n9479.n26 a_n1236_n9479.t15 4.3505
R1234 a_n1236_n9479.n26 a_n1236_n9479.t36 4.3505
R1235 a_n1236_n9479.n27 a_n1236_n9479.t39 4.3505
R1236 a_n1236_n9479.n27 a_n1236_n9479.t3 4.3505
R1237 a_n1236_n9479.n34 a_n1236_n9479.t29 4.3505
R1238 a_n1236_n9479.n34 a_n1236_n9479.t45 4.3505
R1239 a_n1236_n9479.n35 a_n1236_n9479.t40 4.3505
R1240 a_n1236_n9479.n35 a_n1236_n9479.t7 4.3505
R1241 a_n1236_n9479.n69 a_n1236_n9479.t19 4.3505
R1242 a_n1236_n9479.n69 a_n1236_n9479.t44 4.3505
R1243 a_n1236_n9479.n67 a_n1236_n9479.t41 4.3505
R1244 a_n1236_n9479.n67 a_n1236_n9479.t5 4.3505
R1245 a_n1236_n9479.n38 a_n1236_n9479.t21 4.3505
R1246 a_n1236_n9479.n38 a_n1236_n9479.t38 4.3505
R1247 a_n1236_n9479.n39 a_n1236_n9479.t42 4.3505
R1248 a_n1236_n9479.n39 a_n1236_n9479.t1 4.3505
R1249 a_n1236_n9479.n53 a_n1236_n9479.t27 4.3505
R1250 a_n1236_n9479.n53 a_n1236_n9479.t33 4.3505
R1251 a_n1236_n9479.t31 a_n1236_n9479.n84 4.3505
R1252 a_n1236_n9479.n84 a_n1236_n9479.t46 4.3505
R1253 a_n1236_n9479.n9 a_n1236_n9479.n5 2.55258
R1254 a_n1236_n9479.n24 a_n1236_n9479.n14 1.86108
R1255 a_n1236_n9479.n76 a_n1236_n9479.n14 1.86108
R1256 a_n1236_n9479.n76 a_n1236_n9479.n75 1.86108
R1257 a_n1236_n9479.n75 a_n1236_n9479.n15 1.86108
R1258 a_n1236_n9479.n60 a_n1236_n9479.n15 1.86108
R1259 a_n1236_n9479.n60 a_n1236_n9479.n59 1.86108
R1260 a_n1236_n9479.n0 a_n1236_n9479.n9 1.20675
R1261 a_n1236_n9479.n36 a_n1236_n9479.n6 1.0755
R1262 a_n1236_n9479.n12 a_n1236_n9479.n68 1.0755
R1263 a_n1236_n9479.n40 a_n1236_n9479.n10 1.0755
R1264 a_n1236_n9479.n8 a_n1236_n9479.n11 1.0755
R1265 a_n1236_n9479.n2 a_n1236_n9479.n3 1.0755
R1266 a_n1236_n9479.n4 a_n1236_n9479.n1 1.0755
R1267 a_n1236_n9479.n72 a_n1236_n9479.n70 0.759759
R1268 a_n1236_n9479.n74 a_n1236_n9479.n16 0.756673
R1269 a_n1236_n9479.n65 a_n1236_n9479.n37 0.702205
R1270 a_n1236_n9479.n62 a_n1236_n9479.n61 0.700784
R1271 a_n1236_n9479.n80 a_n1236_n9479.n78 0.669534
R1272 a_n1236_n9479.n48 a_n1236_n9479.n46 0.668114
R1273 a_n1236_n9479.n57 a_n1236_n9479.n7 0.666693
R1274 a_n1236_n9479.n82 a_n1236_n9479.n81 0.665273
R1275 a_n1236_n9479.n20 a_n1236_n9479.n19 0.662432
R1276 a_n1236_n9479.n22 a_n1236_n9479.n21 0.661011
R1277 a_n1236_n9479.n56 a_n1236_n9479.n55 0.659208
R1278 a_n1236_n9479.n13 a_n1236_n9479.n74 0.647608
R1279 a_n1236_n9479.n72 a_n1236_n9479.n71 0.645562
R1280 a_n1236_n9479.n23 a_n1236_n9479.n22 0.632599
R1281 a_n1236_n9479.n19 a_n1236_n9479.n18 0.631182
R1282 a_n1236_n9479.n50 a_n1236_n9479.n49 0.629532
R1283 a_n1236_n9479.n82 a_n1236_n9479.n77 0.628338
R1284 a_n1236_n9479.n58 a_n1236_n9479.n7 0.626917
R1285 a_n1236_n9479.n47 a_n1236_n9479.n46 0.625497
R1286 a_n1236_n9479.n79 a_n1236_n9479.n78 0.62408
R1287 a_n1236_n9479.n55 a_n1236_n9479.n42 0.619882
R1288 a_n1236_n9479.n50 a_n1236_n9479.n45 0.594586
R1289 a_n1236_n9479.n63 a_n1236_n9479.n61 0.59283
R1290 a_n1236_n9479.n65 a_n1236_n9479.n64 0.591408
R1291 a_n1236_n9479.n30 a_n1236_n9479.n29 0.580689
R1292 a_n1236_n9479.n33 a_n1236_n9479.n28 0.57833
R1293 a_n1236_n9479.n5 a_n1236_n9479.n4 0.538
R1294 a_n1236_n9479.n6 a_n1236_n9479.n0 0.538
R1295 a_n1236_n9479.n11 a_n1236_n9479.n2 0.537105
R1296 a_n1236_n9479.n1 a_n1236_n9479.n3 0.536664
R1297 a_n1236_n9479.n33 a_n1236_n9479.n32 0.495783
R1298 a_n1236_n9479.n31 a_n1236_n9479.n29 0.493424
R1299 a_n1236_n9479.n71 a_n1236_n9479.n13 0.488952
R1300 a_n1236_n9479.n70 a_n1236_n9479.n16 0.486913
R1301 a_n1236_n9479.n58 a_n1236_n9479.n42 0.476043
R1302 a_n1236_n9479.n57 a_n1236_n9479.n56 0.476043
R1303 a_n1236_n9479.n23 a_n1236_n9479.n18 0.459739
R1304 a_n1236_n9479.n21 a_n1236_n9479.n20 0.459739
R1305 a_n1236_n9479.n79 a_n1236_n9479.n77 0.459739
R1306 a_n1236_n9479.n81 a_n1236_n9479.n80 0.459739
R1307 a_n1236_n9479.n47 a_n1236_n9479.n45 0.459739
R1308 a_n1236_n9479.n49 a_n1236_n9479.n48 0.459739
R1309 a_n1236_n9479.n62 a_n1236_n9479.n37 0.451587
R1310 a_n1236_n9479.n64 a_n1236_n9479.n63 0.451587
R1311 a_n1236_n9479.n54 a_n1236_n9479.n8 0.408833
R1312 a_n1236_n9479.n30 a_n1236_n9479.n28 0.405391
R1313 a_n1236_n9479.n32 a_n1236_n9479.n31 0.405391
R1314 a_n1236_n9479.n73 a_n1236_n9479.n12 0.395292
R1315 a_n1236_n9479.n66 a_n1236_n9479.n10 0.395292
R1316 a_n1236_n9479.n73 a_n1236_n9479.n36 0.143208
R1317 a_n1236_n9479.n68 a_n1236_n9479.n66 0.143208
R1318 3rd_3_OTA_0.vd4.n4 3rd_3_OTA_0.vd4.t4 72.7606
R1319 3rd_3_OTA_0.vd4 3rd_3_OTA_0.vd4.t2 71.6732
R1320 3rd_3_OTA_0.vd4 3rd_3_OTA_0.vd4.n5 62.243
R1321 3rd_3_OTA_0.vd4.n0 3rd_3_OTA_0.vd4.t11 44.7129
R1322 3rd_3_OTA_0.vd4.n0 3rd_3_OTA_0.vd4.t8 44.0566
R1323 3rd_3_OTA_0.vd4.n0 3rd_3_OTA_0.vd4.t12 44.0566
R1324 3rd_3_OTA_0.vd4.n0 3rd_3_OTA_0.vd4.t10 43.8054
R1325 3rd_3_OTA_0.vd4.n1 3rd_3_OTA_0.vd4.t5 19.4751
R1326 3rd_3_OTA_0.vd4.n1 3rd_3_OTA_0.vd4.t6 18.6511
R1327 3rd_3_OTA_0.vd4.n3 3rd_3_OTA_0.vd4.n2 15.6099
R1328 3rd_3_OTA_0.vd4.n5 3rd_3_OTA_0.vd4.t3 11.6005
R1329 3rd_3_OTA_0.vd4.n5 3rd_3_OTA_0.vd4.t1 11.6005
R1330 3rd_3_OTA_0.vd4 3rd_3_OTA_0.vd4.t9 4.23179
R1331 3rd_3_OTA_0.vd4 3rd_3_OTA_0.vd4.n4 2.90758
R1332 3rd_3_OTA_0.vd4 3rd_3_OTA_0.vd4.n0 2.2205
R1333 3rd_3_OTA_0.vd4.n2 3rd_3_OTA_0.vd4.t0 1.90483
R1334 3rd_3_OTA_0.vd4.n2 3rd_3_OTA_0.vd4.t7 1.90483
R1335 3rd_3_OTA_0.vd4.n3 3rd_3_OTA_0.vd4.n1 1.32214
R1336 3rd_3_OTA_0.vd4.n4 3rd_3_OTA_0.vd4.n3 1.28407
R1337 a_7434_1657.n6 a_7434_1657.t12 387.31
R1338 a_7434_1657.n4 a_7434_1657.t5 96.4665
R1339 a_7434_1657.n8 a_7434_1657.t7 96.3265
R1340 a_7434_1657.n0 a_7434_1657.n5 84.9005
R1341 a_7434_1657.n3 a_7434_1657.t2 35.0885
R1342 a_7434_1657.n3 a_7434_1657.t1 34.5018
R1343 a_7434_1657.n9 a_7434_1657.n3 28.9216
R1344 a_7434_1657.n7 a_7434_1657.t6 13.386
R1345 a_7434_1657.n0 a_7434_1657.t10 13.386
R1346 a_7434_1657.n0 a_7434_1657.t8 13.3552
R1347 a_7434_1657.n4 a_7434_1657.t4 13.3552
R1348 a_7434_1657.n5 a_7434_1657.t11 11.4265
R1349 a_7434_1657.n5 a_7434_1657.t9 11.4265
R1350 a_7434_1657.n0 a_7434_1657.n1 2.60415
R1351 a_7434_1657.n9 a_7434_1657.t0 5.8005
R1352 a_7434_1657.t3 a_7434_1657.n9 5.8005
R1353 a_7434_1657.n2 a_7434_1657.n4 5.77814
R1354 a_7434_1657.n7 a_7434_1657.n6 5.54799
R1355 a_7434_1657.n3 a_7434_1657.n0 4.59803
R1356 a_7434_1657.n2 a_7434_1657.n8 3.46037
R1357 a_7434_1657.n6 a_7434_1657.n1 3.00055
R1358 a_7434_1657.n3 a_7434_1657.n2 1.8052
R1359 a_7434_1657.n8 a_7434_1657.n7 1.3961
R1360 a_7434_1657.n1 a_7434_1657.n4 6.41093
R1361 OTA_stage1_0.vd2.t0 OTA_stage1_0.vd2.t2 134.761
R1362 OTA_stage1_0.vd2.t0 OTA_stage1_0.vd2.t1 134.73
R1363 OTA_stage1_0.vd2.t0 OTA_stage1_0.vd2.t5 129.058
R1364 OTA_stage1_0.vd2.t0 OTA_stage1_0.vd2.t3 122.688
R1365 OTA_stage1_0.vd2.t0 OTA_stage1_0.vd2.t6 122.213
R1366 OTA_stage1_0.vd2.t0 OTA_stage1_0.vd2.t4 122.213
R1367 a_n1050_166.n4 a_n1050_166.t10 36.4777
R1368 a_n1050_166.n5 a_n1050_166.t9 35.4327
R1369 a_n1050_166.n4 a_n1050_166.n3 31.3519
R1370 a_n1050_166.n8 a_n1050_166.n7 18.3035
R1371 a_n1050_166.n2 a_n1050_166.n1 18.303
R1372 a_n1050_166.n9 a_n1050_166.n8 17.2098
R1373 a_n1050_166.n2 a_n1050_166.n0 17.208
R1374 a_n1050_166.n6 a_n1050_166.n2 8.938
R1375 a_n1050_166.n3 a_n1050_166.t8 4.08121
R1376 a_n1050_166.n3 a_n1050_166.t0 4.08121
R1377 a_n1050_166.n8 a_n1050_166.n6 3.05142
R1378 a_n1050_166.n6 a_n1050_166.n5 2.2455
R1379 a_n1050_166.n1 a_n1050_166.t2 1.90483
R1380 a_n1050_166.n1 a_n1050_166.t6 1.90483
R1381 a_n1050_166.n0 a_n1050_166.t7 1.90483
R1382 a_n1050_166.n0 a_n1050_166.t4 1.90483
R1383 a_n1050_166.n7 a_n1050_166.t11 1.90483
R1384 a_n1050_166.n7 a_n1050_166.t3 1.90483
R1385 a_n1050_166.t5 a_n1050_166.n9 1.90483
R1386 a_n1050_166.n9 a_n1050_166.t1 1.90483
R1387 a_n1050_166.n5 a_n1050_166.n4 1.0455
R1388 vcc.n213 vcc.n19 17565.9
R1389 vcc.n215 vcc.n19 17565.9
R1390 vcc.n215 vcc.n20 17562.4
R1391 vcc.n213 vcc.n20 17562.4
R1392 vcc.n8 vcc.n5 16027.1
R1393 vcc.n10 vcc.n5 16027.1
R1394 vcc.n8 vcc.n6 16027.1
R1395 vcc.n10 vcc.n6 16027.1
R1396 vcc.n156 vcc.n57 12420
R1397 vcc.n156 vcc.n46 12420
R1398 vcc.n158 vcc.n57 12416.5
R1399 vcc.n158 vcc.n46 12416.5
R1400 vcc.n204 vcc.n34 6349.41
R1401 vcc.n204 vcc.n35 6349.41
R1402 vcc.n202 vcc.n34 6349.41
R1403 vcc.n202 vcc.n35 6349.41
R1404 vcc.n144 vcc.n56 4698.77
R1405 vcc.n94 vcc.n91 3045.88
R1406 vcc.n97 vcc.n91 3045.88
R1407 vcc.n97 vcc.n92 3045.88
R1408 vcc.n135 vcc.n70 2701.93
R1409 vcc.n131 vcc.n72 2372.5
R1410 vcc.n72 vcc.n71 2327.31
R1411 vcc.n103 vcc.n88 2089.41
R1412 vcc.n106 vcc.n87 2089.41
R1413 vcc.n110 vcc.n79 2089.41
R1414 vcc.n113 vcc.n78 2089.41
R1415 vcc.n120 vcc.n119 2089.41
R1416 vcc.n122 vcc.n75 2089.41
R1417 vcc.n177 vcc.n54 2071.76
R1418 vcc.n171 vcc.n162 2071.76
R1419 vcc.n169 vcc.n55 1443.53
R1420 vcc.n169 vcc.n164 1443.53
R1421 vcc.n10 vcc.t21 1353.8
R1422 vcc.t26 vcc.n8 1317.74
R1423 vcc.n9 vcc.t26 1196.03
R1424 vcc.t21 vcc.n9 1159.97
R1425 vcc.n165 vcc.n164 628.236
R1426 vcc.n164 vcc.n54 628.236
R1427 vcc.n171 vcc.n55 628.236
R1428 vcc.n175 vcc.n55 628.236
R1429 vcc.n66 vcc.n65 599.49
R1430 vcc.n7 vcc.n4 415.628
R1431 vcc.n133 vcc.t5 413.37
R1432 vcc.t13 vcc.t15 412.942
R1433 vcc.t17 vcc.t11 412.942
R1434 vcc.n11 vcc.n4 405.284
R1435 vcc.t5 vcc.t32 387.817
R1436 vcc.t15 vcc.n57 319.411
R1437 vcc.t11 vcc.n46 315.507
R1438 vcc.n104 vcc.n87 290.354
R1439 vcc.n105 vcc.n88 290.354
R1440 vcc.n111 vcc.n78 290.354
R1441 vcc.n112 vcc.n79 290.354
R1442 vcc.n122 vcc.n121 290.354
R1443 vcc.n119 vcc.n118 290.354
R1444 vcc.n128 vcc.n127 285.889
R1445 vcc.n132 vcc.n70 268.555
R1446 vcc.n189 vcc.n188 259.036
R1447 vcc.n130 vcc.n129 253.067
R1448 vcc.n129 vcc.n128 248.246
R1449 vcc.n81 vcc.t1 231.379
R1450 vcc.n142 vcc.t49 231.287
R1451 vcc.n61 vcc.t31 231.287
R1452 vcc.n83 vcc.t8 231.287
R1453 vcc.n82 vcc.t37 231.273
R1454 vcc.t35 vcc.t40 216.05
R1455 vcc.t2 vcc.t38 216.05
R1456 vcc.n212 vcc.n16 209.422
R1457 vcc.n157 vcc.t17 208.423
R1458 vcc.n157 vcc.t13 204.519
R1459 vcc.n141 vcc.n62 202.453
R1460 vcc.n7 vcc.n3 183.016
R1461 vcc.n135 vcc.n134 182.202
R1462 vcc.n97 vcc.t0 178.327
R1463 vcc.n12 vcc.n11 176.572
R1464 vcc.t19 vcc.n170 176.514
R1465 vcc.n170 vcc.t45 176.514
R1466 vcc.t40 vcc.n34 174.992
R1467 vcc.t38 vcc.n35 174.992
R1468 vcc.n95 vcc.n94 174.803
R1469 vcc.n177 vcc.n176 173.517
R1470 vcc.n163 vcc.n162 173.517
R1471 vcc.n72 vcc.t9 172.579
R1472 vcc.n173 vcc.n172 166.4
R1473 vcc.n160 vcc.n159 161.126
R1474 vcc.n217 vcc.n17 157.375
R1475 vcc.n168 vcc.n167 153.976
R1476 vcc.n168 vcc.n52 146.825
R1477 vcc.n98 vcc.n90 128.709
R1478 vcc.n166 vcc.n161 124.802
R1479 vcc.n2 vcc.n0 120.891
R1480 vcc.n2 vcc.n1 119.76
R1481 vcc.n130 vcc.n126 118.385
R1482 vcc.n30 vcc.n29 116.722
R1483 vcc.n216 vcc.n18 115.912
R1484 vcc.n99 vcc.n98 115.841
R1485 vcc.n217 vcc.n216 108.909
R1486 vcc.n203 vcc.t35 108.025
R1487 vcc.n203 vcc.t2 108.025
R1488 vcc.n189 vcc.n47 104.57
R1489 vcc.n117 vcc.n73 101.912
R1490 vcc.n51 vcc.t20 98.0045
R1491 vcc.n51 vcc.t46 97.6911
R1492 vcc.n178 vcc.n53 95.9841
R1493 vcc.n25 vcc.n24 87.9664
R1494 vcc.n25 vcc.n18 87.7954
R1495 vcc.n182 vcc.n50 87.2408
R1496 vcc.n185 vcc.n184 87.2408
R1497 vcc.n44 vcc.n43 87.1446
R1498 vcc.n149 vcc.n60 87.1446
R1499 vcc.n160 vcc.n56 85.5143
R1500 vcc.n117 vcc.n116 82.438
R1501 vcc.n108 vcc.n76 73.7015
R1502 vcc.n115 vcc.n76 72.4513
R1503 vcc.n38 vcc.n37 71.8902
R1504 vcc.t29 vcc.n213 71.3347
R1505 vcc.n201 vcc.n36 70.7824
R1506 vcc.n167 vcc.n166 67.0123
R1507 vcc.n167 vcc.n53 67.0123
R1508 vcc.n172 vcc.n161 65.892
R1509 vcc.n208 vcc.n21 65.6211
R1510 vcc.n107 vcc.n80 64.6513
R1511 vcc.n100 vcc.n80 64.1322
R1512 vcc.n128 vcc.n71 61.6672
R1513 vcc.n172 vcc.n171 61.6672
R1514 vcc.n171 vcc.t19 61.6672
R1515 vcc.n54 vcc.n53 61.6672
R1516 vcc.t45 vcc.n54 61.6672
R1517 vcc.n166 vcc.n165 61.6672
R1518 vcc.n175 vcc.n174 61.6672
R1519 vcc.n215 vcc.t25 60.8049
R1520 vcc.n126 vcc.n125 58.2536
R1521 vcc.n146 vcc.n145 57.394
R1522 vcc.n65 vcc.t34 57.1305
R1523 vcc.n65 vcc.t10 57.1305
R1524 vcc.n134 vcc.n71 56.2313
R1525 vcc.n212 vcc.n211 55.3321
R1526 vcc.n176 vcc.n175 54.8697
R1527 vcc.n165 vcc.n163 54.8697
R1528 vcc.t4 vcc.t29 53.6285
R1529 vcc.t25 vcc.t24 53.6285
R1530 vcc.n205 vcc.n33 50.9389
R1531 vcc.n131 vcc.n130 46.2505
R1532 vcc.n93 vcc.n90 45.8455
R1533 vcc.n133 vcc.t9 43.4751
R1534 vcc.n124 vcc.n73 36.2672
R1535 vcc.n155 vcc.n58 35.1478
R1536 vcc.n132 vcc.n131 33.6572
R1537 vcc.n41 vcc.n39 32.1789
R1538 vcc.t24 vcc.n214 32.0794
R1539 vcc.n41 vcc.n40 32.0774
R1540 vcc.n91 vcc.n90 30.8338
R1541 vcc.n96 vcc.n91 30.8338
R1542 vcc.n103 vcc.n102 30.8338
R1543 vcc.n92 vcc.n89 30.8338
R1544 vcc.n75 vcc.n73 30.8338
R1545 vcc.n126 vcc.n70 30.8338
R1546 vcc.n120 vcc.n74 30.8338
R1547 vcc.n114 vcc.n113 30.8338
R1548 vcc.n110 vcc.n109 30.8338
R1549 vcc.n107 vcc.n106 30.8338
R1550 vcc.n30 vcc.n21 30.7043
R1551 vcc.n206 vcc.n205 30.0503
R1552 vcc.n206 vcc.n32 29.6052
R1553 vcc.t32 vcc.n132 29.2303
R1554 vcc.n95 vcc.n92 28.7736
R1555 vcc.n62 vcc.t33 28.5655
R1556 vcc.n62 vcc.t6 28.5655
R1557 vcc.n104 vcc.n103 26.1635
R1558 vcc.n111 vcc.n110 26.1635
R1559 vcc.n113 vcc.n112 26.1635
R1560 vcc.n121 vcc.n120 26.1635
R1561 vcc.n118 vcc.n75 26.1635
R1562 vcc.n106 vcc.n105 26.1635
R1563 vcc.n146 vcc.n144 24.2792
R1564 vcc.n119 vcc.n117 23.1311
R1565 vcc.n87 vcc.n80 23.1255
R1566 vcc.n101 vcc.n88 23.1255
R1567 vcc.n79 vcc.n76 23.1255
R1568 vcc.n123 vcc.n122 23.1255
R1569 vcc.n78 vcc.n77 23.1255
R1570 vcc.n102 vcc.n101 22.5272
R1571 vcc.n214 vcc.t4 21.5497
R1572 vcc.n162 vcc.n161 18.5005
R1573 vcc.n178 vcc.n177 18.5005
R1574 vcc.n169 vcc.n168 18.5005
R1575 vcc.n170 vcc.n169 18.5005
R1576 vcc.n93 vcc.n89 18.4652
R1577 vcc.n179 vcc.n178 18.1802
R1578 vcc.n179 vcc.n52 17.9947
R1579 vcc.n1 vcc.t27 15.8699
R1580 vcc.n1 vcc.t22 15.8699
R1581 vcc.n0 vcc.t28 15.8699
R1582 vcc.n0 vcc.t23 15.8699
R1583 vcc.n137 vcc.n64 14.6377
R1584 vcc.n127 vcc.n69 14.5701
R1585 vcc.n137 vcc.n136 12.7273
R1586 vcc.n125 vcc.n124 12.0598
R1587 vcc.n159 vcc.n48 11.6663
R1588 vcc.n129 vcc.n72 11.563
R1589 vcc.n50 vcc.t47 11.4265
R1590 vcc.n50 vcc.t14 11.4265
R1591 vcc.n184 vcc.t18 11.4265
R1592 vcc.n184 vcc.t42 11.4265
R1593 vcc.n43 vcc.t44 11.4265
R1594 vcc.n43 vcc.t12 11.4265
R1595 vcc.n60 vcc.t16 11.4265
R1596 vcc.n60 vcc.t43 11.4265
R1597 vcc.n98 vcc.n97 10.8829
R1598 vcc.n94 vcc.n93 10.8829
R1599 vcc.n124 vcc.n123 10.3636
R1600 vcc.n11 vcc.n10 10.2783
R1601 vcc.n8 vcc.n7 10.2783
R1602 vcc.n109 vcc.n77 9.97982
R1603 vcc.n123 vcc.n74 9.86377
R1604 vcc.n116 vcc.n115 9.85683
R1605 vcc.n114 vcc.n77 9.83647
R1606 vcc.n134 vcc.n133 9.79085
R1607 vcc.n100 vcc.n99 9.73877
R1608 vcc.n139 vcc.n64 9.6823
R1609 vcc.n108 vcc.n107 9.62493
R1610 vcc.n101 vcc.n86 9.59483
R1611 vcc.n67 vcc 9.58101
R1612 vcc.n29 vcc.n28 9.34567
R1613 vcc.n59 vcc.n58 9.3005
R1614 vcc.n152 vcc.n47 9.3005
R1615 vcc.n49 vcc.n48 9.3005
R1616 vcc.n200 vcc.n199 9.3005
R1617 vcc.n209 vcc.n208 9.3005
R1618 vcc.n26 vcc.n25 9.3005
R1619 vcc.t0 vcc.n96 8.9954
R1620 vcc.n37 vcc.n35 8.04398
R1621 vcc.n36 vcc.n34 8.04398
R1622 vcc.n136 vcc.n135 7.4005
R1623 vcc vcc.n141 7.20708
R1624 vcc.n202 vcc.n201 7.11588
R1625 vcc.n203 vcc.n202 7.11588
R1626 vcc.n205 vcc.n204 7.11588
R1627 vcc.n204 vcc.n203 7.11588
R1628 vcc.n211 vcc.n21 6.56253
R1629 vcc.n174 vcc.n173 5.75273
R1630 vcc.n190 vcc.n46 5.60656
R1631 vcc.n145 vcc.n57 5.60656
R1632 vcc.n24 vcc.n20 5.44168
R1633 vcc.n214 vcc.n20 5.44168
R1634 vcc.n19 vcc.n17 5.44168
R1635 vcc.n214 vcc.n19 5.44168
R1636 vcc.t19 vcc.n163 5.16575
R1637 vcc.n176 vcc.t45 5.16575
R1638 vcc.n201 vcc.n200 4.82369
R1639 vcc.n173 vcc.n160 4.58844
R1640 vcc.n152 vcc.n151 4.5005
R1641 vcc.n183 vcc.n49 4.5005
R1642 vcc.n36 vcc.n33 4.48345
R1643 vcc.n29 vcc.n22 4.42232
R1644 vcc.n105 vcc.t7 4.28573
R1645 vcc.t7 vcc.n104 4.28573
R1646 vcc.n118 vcc.t48 4.28573
R1647 vcc.n121 vcc.t48 4.28573
R1648 vcc.n112 vcc.t30 4.28573
R1649 vcc.t30 vcc.n111 4.28573
R1650 vcc vcc.n143 4.12557
R1651 vcc.n39 vcc.t41 4.08121
R1652 vcc.n39 vcc.t36 4.08121
R1653 vcc.n40 vcc.t3 4.08121
R1654 vcc.n40 vcc.t39 4.08121
R1655 vcc.n194 vcc.n42 3.98496
R1656 vcc.n187 vcc.n45 3.8313
R1657 vcc.n145 vcc.n56 3.22115
R1658 vcc.n180 vcc.n49 3.09113
R1659 vcc.n159 vcc.n158 2.68166
R1660 vcc.n158 vcc.n157 2.68166
R1661 vcc.n156 vcc.n155 2.68166
R1662 vcc.n157 vcc.n156 2.68166
R1663 vcc.n185 vcc.n42 2.55635
R1664 vcc.n200 vcc.n38 1.94833
R1665 vcc.n28 vcc.n27 1.87667
R1666 vcc.n24 vcc.n22 1.86232
R1667 vcc.n193 vcc.n192 1.85463
R1668 vcc.n219 vcc.n218 1.85361
R1669 vcc.n152 vcc.n45 1.78294
R1670 vcc.n96 vcc.n95 1.7705
R1671 vcc.n182 vcc.n181 1.688
R1672 vcc.n213 vcc.n212 1.66717
R1673 vcc.n216 vcc.n215 1.66717
R1674 vcc.n6 vcc.n4 1.63767
R1675 vcc.n9 vcc.n6 1.63767
R1676 vcc.n5 vcc.n3 1.63767
R1677 vcc.n9 vcc.n5 1.63767
R1678 vcc.n85 vcc.n81 1.62503
R1679 vcc.n207 vcc.n206 1.6211
R1680 vcc.n188 vcc.n48 1.45873
R1681 vcc.n15 vcc.n14 1.41806
R1682 vcc.n183 vcc.n182 1.27935
R1683 vcc.n13 vcc 1.27612
R1684 vcc.n221 vcc.n15 1.21641
R1685 vcc.n17 vcc.n16 1.20392
R1686 vcc.n14 vcc.n2 1.20189
R1687 vcc.n37 vcc.n32 1.19816
R1688 vcc.n147 vcc.n59 1.19668
R1689 vcc.n154 vcc.n47 1.19015
R1690 vcc.n147 vcc.n146 1.11733
R1691 vcc.n144 vcc.n58 1.05462
R1692 vcc.n83 vcc.n82 1.00136
R1693 vcc.n210 vcc.n209 0.985286
R1694 vcc.n26 vcc.n23 0.96321
R1695 vcc.n186 vcc.n185 0.963107
R1696 vcc.n174 vcc.n52 0.933293
R1697 vcc.n198 vcc.n197 0.928261
R1698 vcc.n210 vcc.n30 0.875256
R1699 vcc.n211 vcc.n210 0.862026
R1700 vcc.n195 vcc.n194 0.838031
R1701 vcc.n138 vcc.n68 0.813514
R1702 vcc.n153 vcc.n59 0.780009
R1703 vcc.n27 vcc.n26 0.758322
R1704 vcc.n221 vcc.n220 0.680786
R1705 vcc.n136 vcc.n69 0.649348
R1706 vcc.n148 vcc.n147 0.641762
R1707 vcc.n84 vcc.n83 0.612135
R1708 vcc.n190 vcc.n189 0.603552
R1709 vcc.n85 vcc.n84 0.595437
R1710 vcc.n180 vcc.n179 0.58175
R1711 vcc.n196 vcc.n195 0.539263
R1712 vcc.n143 vcc.n61 0.529588
R1713 vcc.n12 vcc.n3 0.492808
R1714 vcc.n197 vcc.n196 0.445398
R1715 vcc.n193 vcc.n44 0.41511
R1716 vcc.n149 vcc.n148 0.407233
R1717 vcc.n84 vcc.n61 0.403016
R1718 vcc.n220 vcc 0.390072
R1719 vcc.n138 vcc.n137 0.358192
R1720 vcc.n150 vcc.n149 0.347903
R1721 vcc.n27 vcc.n18 0.342518
R1722 vcc.n127 vcc.n68 0.332643
R1723 vcc.n195 vcc.n33 0.321789
R1724 vcc.n82 vcc.n81 0.319213
R1725 vcc.n151 vcc.n44 0.314461
R1726 vcc.n155 vcc.n154 0.2565
R1727 vcc.n181 vcc.n180 0.2505
R1728 vcc.n69 vcc.n63 0.239152
R1729 vcc.n125 vcc.n64 0.237537
R1730 vcc.n99 vcc.n89 0.228778
R1731 vcc.n109 vcc.n108 0.212205
R1732 vcc.n143 vcc.n142 0.180531
R1733 vcc.n140 vcc.n63 0.163235
R1734 vcc.n140 vcc.n139 0.1505
R1735 vcc.n68 vcc.n67 0.1505
R1736 vcc.n191 vcc.n190 0.1505
R1737 vcc.n188 vcc.n187 0.148119
R1738 vcc.n208 vcc.n207 0.137839
R1739 vcc.n181 vcc.n51 0.133423
R1740 vcc.n197 vcc.n32 0.129667
R1741 vcc.n23 vcc.n22 0.129667
R1742 vcc.n13 vcc.n12 0.123496
R1743 vcc.n107 vcc.n86 0.114495
R1744 vcc.n66 vcc.n63 0.111978
R1745 vcc.n198 vcc.n38 0.103833
R1746 vcc.n218 vcc.n217 0.0994362
R1747 vcc vcc.n221 0.0953661
R1748 vcc.n219 vcc.n16 0.0866111
R1749 vcc.n115 vcc.n114 0.0831873
R1750 vcc.n102 vcc.n100 0.0819249
R1751 vcc.n86 vcc.n85 0.0678913
R1752 vcc.n192 vcc.n191 0.0666765
R1753 vcc.n187 vcc.n186 0.0638803
R1754 vcc.n142 vcc 0.0571038
R1755 vcc.n67 vcc.n66 0.0519512
R1756 vcc.n116 vcc.n74 0.0501124
R1757 vcc.n199 vcc.n41 0.047375
R1758 vcc.n148 vcc 0.0443375
R1759 vcc.n218 vcc.n15 0.0429528
R1760 vcc.n220 vcc.n219 0.038
R1761 vcc.n139 vcc.n138 0.037915
R1762 vcc.n194 vcc.n193 0.0364015
R1763 vcc.n207 vcc.n31 0.0341957
R1764 vcc.n141 vcc.n140 0.0303556
R1765 vcc.n154 vcc.n153 0.0274565
R1766 vcc.n153 vcc.n152 0.0266936
R1767 vcc.n151 vcc.n150 0.0261494
R1768 vcc.n192 vcc.n42 0.0233659
R1769 vcc.n199 vcc.n198 0.0216694
R1770 vcc.n187 vcc.n49 0.0211422
R1771 vcc.n196 vcc.n31 0.020648
R1772 vcc.n186 vcc.n183 0.0197308
R1773 vcc.n191 vcc.n45 0.0144018
R1774 vcc.n14 vcc.n13 0.0133125
R1775 vcc.n153 vcc.n150 0.0121883
R1776 vcc.n209 vcc.n31 0.00255592
R1777 vcc.n28 vcc.n23 0.00155302
R1778 vin_p.n0 vin_p.t1 21.6012
R1779 vin_p.n0 vin_p.t0 8.85318
R1780 vin_p vin_p.n0 2.55816
R1781 vo3.n0 vo3.t1 98.4603
R1782 vo3.n0 vo3.t2 88.6727
R1783 vo3.n1 vo3.t0 46.53
R1784 vo3.n1 vo3.n0 0.203972
R1785 vo3 vo3.n1 0.107444
R1786 OTA_vref_0.vb1.n1 OTA_vref_0.vb1.n2 71.7516
R1787 OTA_vref_0.vb1.n1 OTA_vref_0.vb1.n3 70.9453
R1788 OTA_vref_0.vb1.n1 OTA_vref_0.vb1.n4 70.9453
R1789 OTA_vref_0.vb1.n0 OTA_vref_0.vb1.t8 68.1062
R1790 OTA_vref_0.vb1.n0 OTA_vref_0.vb1.t9 67.5138
R1791 OTA_vref_0.vb1.n0 OTA_vref_0.vb1.t7 67.5138
R1792 OTA_vref_0.vb1.n0 OTA_vref_0.vb1.t6 67.5138
R1793 OTA_vref_0.vb1.n2 OTA_vref_0.vb1.t5 17.4005
R1794 OTA_vref_0.vb1.n2 OTA_vref_0.vb1.t1 17.4005
R1795 OTA_vref_0.vb1.n3 OTA_vref_0.vb1.t2 17.4005
R1796 OTA_vref_0.vb1.n3 OTA_vref_0.vb1.t0 17.4005
R1797 OTA_vref_0.vb1.n4 OTA_vref_0.vb1.t3 17.4005
R1798 OTA_vref_0.vb1.n4 OTA_vref_0.vb1.t4 17.4005
R1799 OTA_vref_0.vb1 OTA_vref_0.vb1.n0 10.0205
R1800 OTA_vref_0.vb1 OTA_vref_0.vb1.n1 8.74264
R1801 OTA_vref_0.OTA_vref_stage2_0.vr.n4 OTA_vref_0.OTA_vref_stage2_0.vr.t1 651.943
R1802 OTA_vref_0.OTA_vref_stage2_0.vr.n22 OTA_vref_0.OTA_vref_stage2_0.vr.t3 651.74
R1803 OTA_vref_0.OTA_vref_stage2_0.vr.n24 OTA_vref_0.OTA_vref_stage2_0.vr.t23 60.1752
R1804 OTA_vref_0.OTA_vref_stage2_0.vr.n23 OTA_vref_0.OTA_vref_stage2_0.vr.t22 60.1752
R1805 OTA_vref_0.OTA_vref_stage2_0.vr.n14 OTA_vref_0.OTA_vref_stage2_0.vr.t17 28.5589
R1806 OTA_vref_0.OTA_vref_stage2_0.vr.n18 OTA_vref_0.OTA_vref_stage2_0.vr.t7 27.6016
R1807 OTA_vref_0.OTA_vref_stage2_0.vr.n0 OTA_vref_0.OTA_vref_stage2_0.vr.t25 26.8562
R1808 OTA_vref_0.OTA_vref_stage2_0.vr.n0 OTA_vref_0.OTA_vref_stage2_0.vr.t26 26.0492
R1809 OTA_vref_0.OTA_vref_stage2_0.vr.n1 OTA_vref_0.OTA_vref_stage2_0.vr.t21 26.0492
R1810 OTA_vref_0.OTA_vref_stage2_0.vr.n2 OTA_vref_0.OTA_vref_stage2_0.vr.t24 26.0492
R1811 OTA_vref_0.OTA_vref_stage2_0.vr.n3 OTA_vref_0.OTA_vref_stage2_0.vr.t20 26.0492
R1812 OTA_vref_0.OTA_vref_stage2_0.vr.n9 OTA_vref_0.OTA_vref_stage2_0.vr.n8 24.2089
R1813 OTA_vref_0.OTA_vref_stage2_0.vr.n14 OTA_vref_0.OTA_vref_stage2_0.vr.n13 23.2516
R1814 OTA_vref_0.OTA_vref_stage2_0.vr.n15 OTA_vref_0.OTA_vref_stage2_0.vr.n12 23.2516
R1815 OTA_vref_0.OTA_vref_stage2_0.vr.n9 OTA_vref_0.OTA_vref_stage2_0.vr.n7 23.2516
R1816 OTA_vref_0.OTA_vref_stage2_0.vr.n10 OTA_vref_0.OTA_vref_stage2_0.vr.n6 23.2516
R1817 OTA_vref_0.OTA_vref_stage2_0.vr.n11 OTA_vref_0.OTA_vref_stage2_0.vr.n5 23.2516
R1818 OTA_vref_0.OTA_vref_stage2_0.vr.n17 OTA_vref_0.OTA_vref_stage2_0.vr.n16 23.2516
R1819 OTA_vref_0.OTA_vref_stage2_0.vr.n4 OTA_vref_0.OTA_vref_stage2_0.vr.t0 23
R1820 OTA_vref_0.OTA_vref_stage2_0.vr.n21 OTA_vref_0.OTA_vref_stage2_0.vr.t2 23
R1821 OTA_vref_0.OTA_vref_stage2_0.vr.n13 OTA_vref_0.OTA_vref_stage2_0.vr.t10 4.3505
R1822 OTA_vref_0.OTA_vref_stage2_0.vr.n13 OTA_vref_0.OTA_vref_stage2_0.vr.t4 4.3505
R1823 OTA_vref_0.OTA_vref_stage2_0.vr.n12 OTA_vref_0.OTA_vref_stage2_0.vr.t13 4.3505
R1824 OTA_vref_0.OTA_vref_stage2_0.vr.n12 OTA_vref_0.OTA_vref_stage2_0.vr.t18 4.3505
R1825 OTA_vref_0.OTA_vref_stage2_0.vr.n8 OTA_vref_0.OTA_vref_stage2_0.vr.t9 4.3505
R1826 OTA_vref_0.OTA_vref_stage2_0.vr.n8 OTA_vref_0.OTA_vref_stage2_0.vr.t16 4.3505
R1827 OTA_vref_0.OTA_vref_stage2_0.vr.n7 OTA_vref_0.OTA_vref_stage2_0.vr.t8 4.3505
R1828 OTA_vref_0.OTA_vref_stage2_0.vr.n7 OTA_vref_0.OTA_vref_stage2_0.vr.t12 4.3505
R1829 OTA_vref_0.OTA_vref_stage2_0.vr.n6 OTA_vref_0.OTA_vref_stage2_0.vr.t6 4.3505
R1830 OTA_vref_0.OTA_vref_stage2_0.vr.n6 OTA_vref_0.OTA_vref_stage2_0.vr.t14 4.3505
R1831 OTA_vref_0.OTA_vref_stage2_0.vr.n5 OTA_vref_0.OTA_vref_stage2_0.vr.t5 4.3505
R1832 OTA_vref_0.OTA_vref_stage2_0.vr.n5 OTA_vref_0.OTA_vref_stage2_0.vr.t15 4.3505
R1833 OTA_vref_0.OTA_vref_stage2_0.vr.n16 OTA_vref_0.OTA_vref_stage2_0.vr.t11 4.3505
R1834 OTA_vref_0.OTA_vref_stage2_0.vr.n16 OTA_vref_0.OTA_vref_stage2_0.vr.t19 4.3505
R1835 OTA_vref_0.OTA_vref_stage2_0.vr.n20 OTA_vref_0.OTA_vref_stage2_0.vr.n19 3.89276
R1836 OTA_vref_0.OTA_vref_stage2_0.vr.n1 OTA_vref_0.OTA_vref_stage2_0.vr.n0 2.80213
R1837 OTA_vref_0.OTA_vref_stage2_0.vr.n3 OTA_vref_0.OTA_vref_stage2_0.vr.n2 2.76952
R1838 OTA_vref_0.OTA_vref_stage2_0.vr.n2 OTA_vref_0.OTA_vref_stage2_0.vr.n1 2.72333
R1839 OTA_vref_0.OTA_vref_stage2_0.vr.n19 OTA_vref_0.OTA_vref_stage2_0.vr.n11 1.06728
R1840 OTA_vref_0.OTA_vref_stage2_0.vr.n10 OTA_vref_0.OTA_vref_stage2_0.vr.n9 0.957816
R1841 OTA_vref_0.OTA_vref_stage2_0.vr.n11 OTA_vref_0.OTA_vref_stage2_0.vr.n10 0.957816
R1842 OTA_vref_0.OTA_vref_stage2_0.vr.n15 OTA_vref_0.OTA_vref_stage2_0.vr.n14 0.957816
R1843 OTA_vref_0.OTA_vref_stage2_0.vr.n17 OTA_vref_0.OTA_vref_stage2_0.vr.n15 0.957816
R1844 OTA_vref_0.OTA_vref_stage2_0.vr.n18 OTA_vref_0.OTA_vref_stage2_0.vr.n17 0.957816
R1845 OTA_vref_0.OTA_vref_stage2_0.vr.n23 OTA_vref_0.OTA_vref_stage2_0.vr.n22 0.712457
R1846 OTA_vref_0.OTA_vref_stage2_0.vr OTA_vref_0.OTA_vref_stage2_0.vr.n24 0.660826
R1847 OTA_vref_0.OTA_vref_stage2_0.vr OTA_vref_0.OTA_vref_stage2_0.vr.n3 0.617348
R1848 OTA_vref_0.OTA_vref_stage2_0.vr.n19 OTA_vref_0.OTA_vref_stage2_0.vr.n18 0.577487
R1849 OTA_vref_0.OTA_vref_stage2_0.vr.n24 OTA_vref_0.OTA_vref_stage2_0.vr.n23 0.36463
R1850 OTA_vref_0.OTA_vref_stage2_0.vr.n21 OTA_vref_0.OTA_vref_stage2_0.vr.n20 0.240616
R1851 OTA_vref_0.OTA_vref_stage2_0.vr.n20 OTA_vref_0.OTA_vref_stage2_0.vr.n4 0.216527
R1852 OTA_vref_0.OTA_vref_stage2_0.vr.n22 OTA_vref_0.OTA_vref_stage2_0.vr.n21 0.206939
R1853 a_11275_n2439.t0 a_11275_n2439.t1 50.1091
R1854 3rd_3_OTA_0.vd1.n0 3rd_3_OTA_0.vd1.t0 138.714
R1855 3rd_3_OTA_0.vd1.n1 3rd_3_OTA_0.vd1.t1 136.073
R1856 3rd_3_OTA_0.vd1.n1 3rd_3_OTA_0.vd1.t6 122.216
R1857 3rd_3_OTA_0.vd1.n1 3rd_3_OTA_0.vd1.t4 122.216
R1858 3rd_3_OTA_0.vd1.n1 3rd_3_OTA_0.vd1.t5 121.828
R1859 3rd_3_OTA_0.vd1.n1 3rd_3_OTA_0.vd1.t7 121.828
R1860 3rd_3_OTA_0.vd1.n0 3rd_3_OTA_0.vd1.t3 19.5045
R1861 3rd_3_OTA_0.vd1.n1 3rd_3_OTA_0.vd1.t2 17.559
R1862 3rd_3_OTA_0.vd1.n1 3rd_3_OTA_0.vd1.n0 11.1867
R1863 3rd_3_OTA_0.vd1 3rd_3_OTA_0.vd1.n1 9.24116
R1864 vin_n.n0 vin_n.t1 21.0692
R1865 vin_n.n0 vin_n.t0 8.85313
R1866 vin_n vin_n.n0 2.40005
C0 a_2382_n6868# a_2470_n7958# 0.097592f
C1 a_2382_n4288# vcc 0.368035f
C2 a_2382_n5578# a_2382_n6868# 0.154516f
C3 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage2_0.vr 9.256969f
C4 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vr 2.20674f
C5 a_2470_n5378# OTA_vref_0.vb1 0.038035f
C6 a_11847_n1701# vcc 0.836592f
C7 OTA_vref_0.OTA_vref_stage2_0.vr 3rd_3_OTA_0.vd3 0.001587f
C8 a_9040_n3397# 3rd_3_OTA_0.vd4 1.93202f
C9 vin_n 3rd_3_OTA_0.vd1 0.784618f
C10 a_2470_n7958# OTA_vref_0.OTA_vref_stage2_0.vr 0.008049f
C11 a_2382_n5578# OTA_vref_0.OTA_vref_stage2_0.vr 0.334808f
C12 a_2382_n6868# vcc 0.318981f
C13 vin_n 3rd_3_OTA_0.vb 0.605449f
C14 vin_p vin_n 2.36446f
C15 a_9040_n3397# 3rd_3_OTA_0.vd1 0.006984f
C16 3rd_3_OTA_0.vd3 3rd_3_OTA_0.vd4 9.51896f
C17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 3rd_3_OTA_0.vb 0.006315f
C18 a_2382_n4288# OTA_vref_0.OTA_vref_stage2_0.vr 0.368863f
C19 OTA_vref_0.OTA_vref_stage2_0.vref0 3rd_3_OTA_0.vb 4.32e-19
C20 a_9040_n3397# 3rd_3_OTA_0.vb 1.48336f
C21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2382_n8158# 0.032619f
C22 a_2382_n8158# OTA_vref_0.OTA_vref_stage2_0.vref0 0.112341f
C23 3rd_3_OTA_0.vd3 3rd_3_OTA_0.vd1 1.22886f
C24 3rd_3_OTA_0.vd1 vo3 0.366634f
C25 a_n10077_1624# 3rd_3_OTA_0.vd1 0.118468f
C26 vcc OTA_vref_0.OTA_vref_stage2_0.vr 11.398701f
C27 3rd_3_OTA_0.vd3 3rd_3_OTA_0.vb 0.483395f
C28 a_2382_n4288# 3rd_3_OTA_0.vd4 2.1e-20
C29 a_n10077_1624# 3rd_3_OTA_0.vb 0.443825f
C30 a_2470_n5378# OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 6.62e-20
C31 a_2470_n5378# OTA_vref_0.OTA_vref_stage2_0.vref0 0.00151f
C32 vin_p a_n10077_1624# 1.68092f
C33 a_2470_n7958# a_2382_n8158# 1.53765f
C34 a_11847_n1701# 3rd_3_OTA_0.vd4 1.15e-20
C35 a_2382_n5578# 3rd_3_OTA_0.vb 3.04e-19
C36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.vb1 6.15e-19
C37 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.vb1 0.006422f
C38 a_2382_n6868# OTA_vref_0.OTA_vref_stage2_0.vr 0.341152f
C39 vcc 3rd_3_OTA_0.vd4 4.40467f
C40 a_2382_n4288# 3rd_3_OTA_0.vb 1.67298f
C41 a_11847_n1701# 3rd_3_OTA_0.vd1 0.011993f
C42 OTA_vref_0.vb1 3rd_3_OTA_0.vd3 0.316815f
C43 a_2470_n5378# a_2382_n5578# 1.53005f
C44 a_2470_n7958# OTA_vref_0.vb1 0.056235f
C45 vcc 3rd_3_OTA_0.vd1 8.20565f
C46 a_2382_n5578# OTA_vref_0.vb1 0.106848f
C47 vcc 3rd_3_OTA_0.vb 0.434712f
C48 vcc a_2382_n8158# 0.3278f
C49 vin_p vcc 0.018752f
C50 a_2382_n4288# a_2470_n5378# 0.10061f
C51 a_2382_n6868# a_2382_n8158# 0.154705f
C52 a_2470_n5378# vcc 0.034455f
C53 vcc OTA_vref_0.vb1 8.322209f
C54 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage2_0.vref0 16.2573f
C55 a_2470_n5378# a_2382_n6868# 1.04e-19
C56 vin_n a_n10077_1624# 1.47482f
C57 a_2382_n6868# OTA_vref_0.vb1 1.61373f
C58 OTA_vref_0.OTA_vref_stage2_0.vr 3rd_3_OTA_0.vb 0.233485f
C59 a_2382_n8158# OTA_vref_0.OTA_vref_stage2_0.vr 0.33605f
C60 a_9040_n3397# 3rd_3_OTA_0.vd3 1.97254f
C61 a_9040_n3397# vo3 0.004168f
C62 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_2470_n7958# 0.003419f
C63 a_2470_n7958# OTA_vref_0.OTA_vref_stage2_0.vref0 0.037994f
C64 a_2382_n5578# OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.007176f
C65 a_2382_n5578# OTA_vref_0.OTA_vref_stage2_0.vref0 0.011315f
C66 3rd_3_OTA_0.vd4 3rd_3_OTA_0.vd1 15.7657f
C67 3rd_3_OTA_0.vd4 3rd_3_OTA_0.vb 0.322891f
C68 a_2470_n5378# OTA_vref_0.OTA_vref_stage2_0.vr 0.008037f
C69 a_2382_n4288# OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.002329f
C70 OTA_vref_0.OTA_vref_stage2_0.vr OTA_vref_0.vb1 0.062593f
C71 vin_n vcc 0.018448f
C72 a_9040_n3397# a_11847_n1701# 0.016974f
C73 3rd_3_OTA_0.vb 3rd_3_OTA_0.vd1 0.237308f
C74 vin_p 3rd_3_OTA_0.vd1 0.13787f
C75 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter vcc 0.512021f
C76 a_9040_n3397# vcc 0.101608f
C77 vcc OTA_vref_0.OTA_vref_stage2_0.vref0 0.030224f
C78 a_2382_n4288# 3rd_3_OTA_0.vd3 0.00236f
C79 vin_p 3rd_3_OTA_0.vb 0.39332f
C80 OTA_vref_0.vb1 3rd_3_OTA_0.vd4 0.226739f
C81 a_11847_n1701# 3rd_3_OTA_0.vd3 1.12e-19
C82 a_11847_n1701# vo3 0.159655f
C83 a_2382_n4288# a_2382_n5578# 0.154422f
C84 a_2382_n6868# OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.009524f
C85 a_2382_n6868# OTA_vref_0.OTA_vref_stage2_0.vref0 0.010991f
C86 vcc 3rd_3_OTA_0.vd3 4.62835f
C87 vcc vo3 0.594996f
C88 vcc a_n10077_1624# 5.64e-19
C89 a_2470_n5378# 3rd_3_OTA_0.vb 0.036384f
C90 vcc a_2470_n7958# 0.034292f
C91 a_2382_n5578# vcc 0.335707f
C92 OTA_vref_0.vb1 3rd_3_OTA_0.vb 0.111837f
C93 a_2382_n8158# OTA_vref_0.vb1 0.034229f
C94 vo3 vss 2.83219f
C95 vin_n vss 15.210062f
C96 vin_p vss 14.908583f
C97 vcc vss 0.225p
C98 a_2382_n8158# vss 3.83372f
C99 a_2470_n7958# vss 0.471548f
C100 a_2382_n6868# vss 3.70817f
C101 a_2382_n5578# vss 3.70757f
C102 a_2470_n5378# vss 0.471213f
C103 a_2382_n4288# vss 3.74312f
C104 OTA_vref_0.OTA_vref_stage2_0.vref0 vss 11.528516f
C105 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter vss 25.278364f
C106 OTA_vref_0.OTA_vref_stage2_0.vr vss 12.014772f
C107 a_11847_n1701# vss 1.4749f
C108 a_9040_n3397# vss 5.41946f
C109 OTA_vref_0.vb1 vss 8.843204f
C110 3rd_3_OTA_0.vd3 vss 48.684086f
C111 3rd_3_OTA_0.vd4 vss 19.921677f
C112 3rd_3_OTA_0.vb vss 18.068f
C113 a_n10077_1624# vss 3.49104f
C114 3rd_3_OTA_0.vd1 vss 63.1497f
C115 vin_n.t1 vss 0.869123f
C116 vin_n.t0 vss 0.457268f
C117 vin_n.n0 vss 1.00705f
C118 3rd_3_OTA_0.vd1.n0 vss 1.9415f
C119 3rd_3_OTA_0.vd1.n1 vss 19.1674f
C120 3rd_3_OTA_0.vd1.t1 vss 0.043314f
C121 3rd_3_OTA_0.vd1.t0 vss 0.047902f
C122 3rd_3_OTA_0.vd1.t3 vss 0.356063f
C123 3rd_3_OTA_0.vd1.t2 vss 0.217646f
C124 3rd_3_OTA_0.vd1.t5 vss 1.58819f
C125 3rd_3_OTA_0.vd1.t6 vss 1.59871f
C126 3rd_3_OTA_0.vd1.t4 vss 1.59871f
C127 3rd_3_OTA_0.vd1.t7 vss 1.58819f
C128 a_11275_n2439.t1 vss 26.271801f
C129 a_11275_n2439.t0 vss 0.028206f
C130 OTA_vref_0.OTA_vref_stage2_0.vr.t25 vss 0.60782f
C131 OTA_vref_0.OTA_vref_stage2_0.vr.t26 vss 0.584499f
C132 OTA_vref_0.OTA_vref_stage2_0.vr.n0 vss 1.65263f
C133 OTA_vref_0.OTA_vref_stage2_0.vr.t21 vss 0.584499f
C134 OTA_vref_0.OTA_vref_stage2_0.vr.n1 vss 0.976322f
C135 OTA_vref_0.OTA_vref_stage2_0.vr.t24 vss 0.584499f
C136 OTA_vref_0.OTA_vref_stage2_0.vr.n2 vss 0.97502f
C137 OTA_vref_0.OTA_vref_stage2_0.vr.t20 vss 0.584499f
C138 OTA_vref_0.OTA_vref_stage2_0.vr.n3 vss 0.890892f
C139 OTA_vref_0.OTA_vref_stage2_0.vr.t23 vss 0.303436f
C140 OTA_vref_0.OTA_vref_stage2_0.vr.t22 vss 0.303436f
C141 OTA_vref_0.OTA_vref_stage2_0.vr.t3 vss 0.025841f
C142 OTA_vref_0.OTA_vref_stage2_0.vr.t2 vss 0.458739f
C143 OTA_vref_0.OTA_vref_stage2_0.vr.t0 vss 0.458739f
C144 OTA_vref_0.OTA_vref_stage2_0.vr.t1 vss 0.02587f
C145 OTA_vref_0.OTA_vref_stage2_0.vr.n4 vss 0.832695f
C146 OTA_vref_0.OTA_vref_stage2_0.vr.t5 vss 0.054748f
C147 OTA_vref_0.OTA_vref_stage2_0.vr.t15 vss 0.054748f
C148 OTA_vref_0.OTA_vref_stage2_0.vr.n5 vss 0.20797f
C149 OTA_vref_0.OTA_vref_stage2_0.vr.t6 vss 0.054748f
C150 OTA_vref_0.OTA_vref_stage2_0.vr.t14 vss 0.054748f
C151 OTA_vref_0.OTA_vref_stage2_0.vr.n6 vss 0.20797f
C152 OTA_vref_0.OTA_vref_stage2_0.vr.t8 vss 0.054748f
C153 OTA_vref_0.OTA_vref_stage2_0.vr.t12 vss 0.054748f
C154 OTA_vref_0.OTA_vref_stage2_0.vr.n7 vss 0.20797f
C155 OTA_vref_0.OTA_vref_stage2_0.vr.t9 vss 0.054748f
C156 OTA_vref_0.OTA_vref_stage2_0.vr.t16 vss 0.054748f
C157 OTA_vref_0.OTA_vref_stage2_0.vr.n8 vss 0.236203f
C158 OTA_vref_0.OTA_vref_stage2_0.vr.n9 vss 1.66546f
C159 OTA_vref_0.OTA_vref_stage2_0.vr.n10 vss 0.97974f
C160 OTA_vref_0.OTA_vref_stage2_0.vr.n11 vss 1.0171f
C161 OTA_vref_0.OTA_vref_stage2_0.vr.t7 vss 0.276061f
C162 OTA_vref_0.OTA_vref_stage2_0.vr.t13 vss 0.054748f
C163 OTA_vref_0.OTA_vref_stage2_0.vr.t18 vss 0.054748f
C164 OTA_vref_0.OTA_vref_stage2_0.vr.n12 vss 0.20797f
C165 OTA_vref_0.OTA_vref_stage2_0.vr.t10 vss 0.054748f
C166 OTA_vref_0.OTA_vref_stage2_0.vr.t4 vss 0.054748f
C167 OTA_vref_0.OTA_vref_stage2_0.vr.n13 vss 0.20797f
C168 OTA_vref_0.OTA_vref_stage2_0.vr.t17 vss 0.301381f
C169 OTA_vref_0.OTA_vref_stage2_0.vr.n14 vss 1.70977f
C170 OTA_vref_0.OTA_vref_stage2_0.vr.n15 vss 0.97974f
C171 OTA_vref_0.OTA_vref_stage2_0.vr.t11 vss 0.054748f
C172 OTA_vref_0.OTA_vref_stage2_0.vr.t19 vss 0.054748f
C173 OTA_vref_0.OTA_vref_stage2_0.vr.n16 vss 0.20797f
C174 OTA_vref_0.OTA_vref_stage2_0.vr.n17 vss 0.97974f
C175 OTA_vref_0.OTA_vref_stage2_0.vr.n18 vss 0.920416f
C176 OTA_vref_0.OTA_vref_stage2_0.vr.n19 vss 1.68401f
C177 OTA_vref_0.OTA_vref_stage2_0.vr.n20 vss 0.843703f
C178 OTA_vref_0.OTA_vref_stage2_0.vr.n21 vss 0.768139f
C179 OTA_vref_0.OTA_vref_stage2_0.vr.n22 vss 0.122166f
C180 OTA_vref_0.OTA_vref_stage2_0.vr.n23 vss 0.367868f
C181 OTA_vref_0.OTA_vref_stage2_0.vr.n24 vss 0.365806f
C182 OTA_vref_0.vb1.n0 vss 5.75346f
C183 OTA_vref_0.vb1.n1 vss 0.352136f
C184 OTA_vref_0.vb1.t8 vss 0.858318f
C185 OTA_vref_0.vb1.t9 vss 0.846486f
C186 OTA_vref_0.vb1.t7 vss 0.846486f
C187 OTA_vref_0.vb1.t6 vss 0.846486f
C188 OTA_vref_0.vb1.t5 vss 0.007035f
C189 OTA_vref_0.vb1.t1 vss 0.007035f
C190 OTA_vref_0.vb1.n2 vss 0.018857f
C191 OTA_vref_0.vb1.t2 vss 0.007035f
C192 OTA_vref_0.vb1.t0 vss 0.007035f
C193 OTA_vref_0.vb1.n3 vss 0.017824f
C194 OTA_vref_0.vb1.t3 vss 0.007035f
C195 OTA_vref_0.vb1.t4 vss 0.007035f
C196 OTA_vref_0.vb1.n4 vss 0.017824f
C197 vin_p.t1 vss 0.872831f
C198 vin_p.t0 vss 0.458725f
C199 vin_p.n0 vss 1.00306f
C200 vcc.t28 vss 0.00408f
C201 vcc.t23 vss 0.00408f
C202 vcc.n0 vss 0.008952f
C203 vcc.t27 vss 0.00408f
C204 vcc.t22 vss 0.00408f
C205 vcc.n1 vss 0.008524f
C206 vcc.n2 vss 0.094597f
C207 vcc.n3 vss 0.632551f
C208 vcc.n4 vss 0.453591f
C209 vcc.n5 vss 0.120795f
C210 vcc.n6 vss 0.120795f
C211 vcc.n7 vss 0.83274f
C212 vcc.n8 vss 1.43449f
C213 vcc.t26 vss 2.25072f
C214 vcc.n9 vss 2.10841f
C215 vcc.t21 vss 2.25043f
C216 vcc.n10 vss 1.43248f
C217 vcc.n11 vss 0.89715f
C218 vcc.n12 vss 0.80164f
C219 vcc.n13 vss 1.07672f
C220 vcc.n14 vss 0.726614f
C221 vcc.n15 vss 0.661059f
C222 vcc.n16 vss 0.419212f
C223 vcc.n17 vss 0.277623f
C224 vcc.n18 vss 0.741935f
C225 vcc.n19 vss 0.132939f
C226 vcc.n20 vss 0.132912f
C227 vcc.n21 vss 0.606179f
C228 vcc.n22 vss 0.005222f
C229 vcc.n23 vss 0.077426f
C230 vcc.n24 vss 0.075659f
C231 vcc.n25 vss 0.241686f
C232 vcc.n26 vss 0.189623f
C233 vcc.n27 vss 0.285709f
C234 vcc.n28 vss 0.474937f
C235 vcc.n29 vss 0.143822f
C236 vcc.n30 vss 0.478605f
C237 vcc.n31 vss 0.006415f
C238 vcc.n32 vss 0.109988f
C239 vcc.n33 vss 0.856411f
C240 vcc.n34 vss 0.342239f
C241 vcc.n35 vss 0.342239f
C242 vcc.t40 vss 0.546372f
C243 vcc.t35 vss 0.450331f
C244 vcc.n36 vss 0.372929f
C245 vcc.n37 vss 0.256975f
C246 vcc.n38 vss 0.212378f
C247 vcc.t41 vss 0.015865f
C248 vcc.t36 vss 0.015865f
C249 vcc.n39 vss 0.041211f
C250 vcc.t3 vss 0.015865f
C251 vcc.t39 vss 0.015865f
C252 vcc.n40 vss 0.040451f
C253 vcc.n41 vss 0.64728f
C254 vcc.n42 vss 0.127946f
C255 vcc.t44 vss 0.005666f
C256 vcc.t12 vss 0.005666f
C257 vcc.n43 vss 0.01228f
C258 vcc.n44 vss 0.383059f
C259 vcc.n45 vss 0.365549f
C260 vcc.n46 vss 0.964808f
C261 vcc.n47 vss 1.46047f
C262 vcc.n48 vss 0.010002f
C263 vcc.n49 vss 0.118031f
C264 vcc.t47 vss 0.005666f
C265 vcc.t14 vss 0.005666f
C266 vcc.n50 vss 0.01233f
C267 vcc.t20 vss 0.022588f
C268 vcc.t46 vss 0.022407f
C269 vcc.n51 vss 0.118431f
C270 vcc.n52 vss 0.022593f
C271 vcc.n53 vss 0.016411f
C272 vcc.n54 vss 0.010479f
C273 vcc.t45 vss 0.143356f
C274 vcc.n55 vss 0.010164f
C275 vcc.n56 vss 0.069257f
C276 vcc.n57 vss 0.944443f
C277 vcc.t15 vss 1.78619f
C278 vcc.t13 vss 1.50469f
C279 vcc.t11 vss 1.77724f
C280 vcc.t17 vss 1.5142f
C281 vcc.n58 vss 0.798495f
C282 vcc.n59 vss 0.388785f
C283 vcc.t16 vss 0.005666f
C284 vcc.t43 vss 0.005666f
C285 vcc.n60 vss 0.01228f
C286 vcc.t31 vss 0.008497f
C287 vcc.n61 vss 0.099887f
C288 vcc.t49 vss 0.008497f
C289 vcc.t33 vss 0.002266f
C290 vcc.t6 vss 0.002266f
C291 vcc.n62 vss 0.004835f
C292 vcc.n63 vss 0.298189f
C293 vcc.n64 vss 0.085716f
C294 vcc.t34 vss 0.001133f
C295 vcc.t10 vss 0.001133f
C296 vcc.n65 vss 0.002374f
C297 vcc.n66 vss 0.092952f
C298 vcc.n67 vss 0.16816f
C299 vcc.n68 vss 0.110389f
C300 vcc.n69 vss 0.163684f
C301 vcc.n70 vss 0.111178f
C302 vcc.n71 vss 0.044206f
C303 vcc.t9 vss 0.127156f
C304 vcc.n72 vss 0.175966f
C305 vcc.n73 vss 0.025384f
C306 vcc.n74 vss 0.069822f
C307 vcc.n75 vss 0.016228f
C308 vcc.t48 vss 0.180208f
C309 vcc.n76 vss 0.027477f
C310 vcc.n77 vss 0.109526f
C311 vcc.n78 vss 0.123486f
C312 vcc.n79 vss 0.123486f
C313 vcc.n80 vss 0.029378f
C314 vcc.t1 vss 0.008544f
C315 vcc.n81 vss 0.322107f
C316 vcc.t8 vss 0.008497f
C317 vcc.t37 vss 0.008496f
C318 vcc.n82 vss 0.138361f
C319 vcc.n83 vss 0.154083f
C320 vcc.n84 vss 0.31963f
C321 vcc.n85 vss 0.177111f
C322 vcc.n86 vss 0.071348f
C323 vcc.n87 vss 0.123486f
C324 vcc.n88 vss 0.123486f
C325 vcc.n89 vss 0.119222f
C326 vcc.n90 vss 0.099146f
C327 vcc.n91 vss 0.023568f
C328 vcc.n92 vss 0.023568f
C329 vcc.n93 vss 0.283597f
C330 vcc.n94 vss 0.216749f
C331 vcc.n96 vss 0.155726f
C332 vcc.t0 vss 0.148731f
C333 vcc.n97 vss 0.206576f
C334 vcc.n98 vss 0.049158f
C335 vcc.n99 vss 0.212076f
C336 vcc.n100 vss 0.203122f
C337 vcc.n101 vss 0.132996f
C338 vcc.n102 vss 0.047617f
C339 vcc.n103 vss 0.016228f
C340 vcc.t7 vss 0.180208f
C341 vcc.n106 vss 0.016228f
C342 vcc.n107 vss 0.200703f
C343 vcc.n108 vss 0.200898f
C344 vcc.n109 vss 0.070263f
C345 vcc.n110 vss 0.016228f
C346 vcc.t30 vss 0.180208f
C347 vcc.n113 vss 0.016228f
C348 vcc.n114 vss 0.07107f
C349 vcc.n115 vss 0.197766f
C350 vcc.n116 vss 0.196159f
C351 vcc.n117 vss 0.028744f
C352 vcc.n119 vss 0.123488f
C353 vcc.n120 vss 0.016228f
C354 vcc.n122 vss 0.123486f
C355 vcc.n123 vss 0.111496f
C356 vcc.n124 vss 0.132775f
C357 vcc.n125 vss 0.074326f
C358 vcc.n126 vss 0.013291f
C359 vcc.n127 vss 0.265016f
C360 vcc.n128 vss 0.031885f
C361 vcc.n129 vss 0.035717f
C362 vcc.n130 vss 0.026735f
C363 vcc.n131 vss 0.026735f
C364 vcc.n132 vss 0.040538f
C365 vcc.t32 vss 0.091833f
C366 vcc.t5 vss 0.131633f
C367 vcc.n133 vss 0.144988f
C368 vcc.n134 vss 0.06902f
C369 vcc.n135 vss 0.216205f
C370 vcc.n136 vss 0.076653f
C371 vcc.n137 vss 0.155432f
C372 vcc.n138 vss 0.056853f
C373 vcc.n139 vss 0.059273f
C374 vcc.n140 vss 0.087396f
C375 vcc.n141 vss 0.156454f
C376 vcc.n142 vss 0.044963f
C377 vcc.n143 vss 4.31925f
C378 vcc.n144 vss 0.094328f
C379 vcc.n145 vss 0.044457f
C380 vcc.n146 vss 0.084927f
C381 vcc.n147 vss 0.077964f
C382 vcc.n148 vss 0.277823f
C383 vcc.n149 vss 0.394534f
C384 vcc.n150 vss 0.172862f
C385 vcc.n151 vss 0.157365f
C386 vcc.n152 vss 0.596784f
C387 vcc.n153 vss 0.357986f
C388 vcc.n154 vss 0.031887f
C389 vcc.n155 vss 0.780891f
C390 vcc.n156 vss 0.093799f
C391 vcc.n157 vss 1.00629f
C392 vcc.n158 vss 0.093772f
C393 vcc.n159 vss 0.131745f
C394 vcc.n160 vss 0.248316f
C395 vcc.n161 vss 0.040138f
C396 vcc.n162 vss 0.112103f
C397 vcc.n164 vss 0.010164f
C398 vcc.n165 vss 0.010479f
C399 vcc.n166 vss 0.01371f
C400 vcc.n167 vss 0.010164f
C401 vcc.n168 vss 0.010616f
C402 vcc.n169 vss 0.010868f
C403 vcc.n170 vss 0.133271f
C404 vcc.t19 vss 0.143356f
C405 vcc.n171 vss 0.010479f
C406 vcc.n172 vss 0.140585f
C407 vcc.n173 vss 0.079819f
C408 vcc.n174 vss 0.049804f
C409 vcc.n175 vss 0.010479f
C410 vcc.n177 vss 0.112103f
C411 vcc.n178 vss 0.050768f
C412 vcc.n179 vss 0.021031f
C413 vcc.n180 vss 0.186334f
C414 vcc.n181 vss 0.039044f
C415 vcc.n182 vss 0.173334f
C416 vcc.n183 vss 0.055549f
C417 vcc.t18 vss 0.005666f
C418 vcc.t42 vss 0.005666f
C419 vcc.n184 vss 0.01233f
C420 vcc.n185 vss 0.199477f
C421 vcc.n186 vss 0.042016f
C422 vcc.n187 vss 0.143622f
C423 vcc.n188 vss 0.204977f
C424 vcc.n189 vss 0.558152f
C425 vcc.n190 vss 0.071614f
C426 vcc.n191 vss 0.046695f
C427 vcc.n192 vss 0.039956f
C428 vcc.n193 vss 0.247267f
C429 vcc.n194 vss 0.490484f
C430 vcc.n195 vss 1.31065f
C431 vcc.n196 vss 0.693266f
C432 vcc.n197 vss 0.270645f
C433 vcc.n198 vss 0.192437f
C434 vcc.n199 vss 0.206419f
C435 vcc.n200 vss 0.015746f
C436 vcc.n201 vss 0.232814f
C437 vcc.n202 vss 0.04823f
C438 vcc.t38 vss 0.546372f
C439 vcc.t2 vss 0.450331f
C440 vcc.n203 vss 0.300221f
C441 vcc.n204 vss 0.04823f
C442 vcc.n205 vss 0.560855f
C443 vcc.n206 vss 0.31567f
C444 vcc.n207 vss 0.011654f
C445 vcc.n208 vss 0.435942f
C446 vcc.n209 vss 0.285104f
C447 vcc.n210 vss 0.437443f
C448 vcc.n211 vss 0.199221f
C449 vcc.n212 vss 0.60234f
C450 vcc.n213 vss 2.62868f
C451 vcc.t29 vss 3.11291f
C452 vcc.t4 vss 1.86163f
C453 vcc.n214 vss 1.328f
C454 vcc.t24 vss 2.12238f
C455 vcc.t25 vss 2.85087f
C456 vcc.n215 vss 2.2055f
C457 vcc.n216 vss 0.375817f
C458 vcc.n217 vss 0.453986f
C459 vcc.n218 vss 0.459081f
C460 vcc.n219 vss 0.470702f
C461 vcc.n220 vss 0.767997f
C462 vcc.n221 vss 0.224247f
C463 a_n1050_166.t1 vss 0.216942f
C464 a_n1050_166.t7 vss 0.216942f
C465 a_n1050_166.t4 vss 0.216942f
C466 a_n1050_166.n0 vss 0.671366f
C467 a_n1050_166.t2 vss 0.216942f
C468 a_n1050_166.t6 vss 0.216942f
C469 a_n1050_166.n1 vss 0.762068f
C470 a_n1050_166.n2 vss 4.7253f
C471 a_n1050_166.t9 vss 0.399519f
C472 a_n1050_166.t8 vss 0.10124f
C473 a_n1050_166.t0 vss 0.10124f
C474 a_n1050_166.n3 vss 0.235864f
C475 a_n1050_166.t10 vss 0.427351f
C476 a_n1050_166.n4 vss 2.07187f
C477 a_n1050_166.n5 vss 1.4064f
C478 a_n1050_166.n6 vss 2.8881f
C479 a_n1050_166.t11 vss 0.216942f
C480 a_n1050_166.t3 vss 0.216942f
C481 a_n1050_166.n7 vss 0.76209f
C482 a_n1050_166.n8 vss 3.54056f
C483 a_n1050_166.n9 vss 0.671495f
C484 a_n1050_166.t5 vss 0.216942f
C485 OTA_stage1_0.vd2.t0 vss 38.949104f
C486 OTA_stage1_0.vd2.t3 vss 1.328f
C487 OTA_stage1_0.vd2.t4 vss 1.32133f
C488 OTA_stage1_0.vd2.t6 vss 1.32133f
C489 OTA_stage1_0.vd2.t5 vss 1.31275f
C490 OTA_stage1_0.vd2.t2 vss 0.033752f
C491 OTA_stage1_0.vd2.t1 vss 0.03374f
C492 a_7434_1657.n0 vss 4.28231f
C493 a_7434_1657.n1 vss 0.749832f
C494 a_7434_1657.n2 vss 1.31373f
C495 a_7434_1657.n3 vss 3.19052f
C496 a_7434_1657.n4 vss 2.45343f
C497 a_7434_1657.t0 vss 0.022035f
C498 a_7434_1657.t5 vss 0.067647f
C499 a_7434_1657.t12 vss 0.104031f
C500 a_7434_1657.t4 vss 1.21697f
C501 a_7434_1657.t10 vss 1.2203f
C502 a_7434_1657.t11 vss 0.018363f
C503 a_7434_1657.t9 vss 0.018363f
C504 a_7434_1657.n5 vss 0.03741f
C505 a_7434_1657.t8 vss 1.21697f
C506 a_7434_1657.n6 vss 0.977679f
C507 a_7434_1657.t6 vss 1.22017f
C508 a_7434_1657.n7 vss 1.98638f
C509 a_7434_1657.t7 vss 0.06752f
C510 a_7434_1657.n8 vss 0.144523f
C511 a_7434_1657.t2 vss 0.106961f
C512 a_7434_1657.t1 vss 0.098082f
C513 a_7434_1657.n9 vss 0.064739f
C514 a_7434_1657.t3 vss 0.022035f
C515 3rd_3_OTA_0.vd4.n0 vss 2.57228f
C516 3rd_3_OTA_0.vd4.t11 vss 0.527637f
C517 3rd_3_OTA_0.vd4.t12 vss 0.524989f
C518 3rd_3_OTA_0.vd4.t8 vss 0.52535f
C519 3rd_3_OTA_0.vd4.t10 vss 0.51535f
C520 3rd_3_OTA_0.vd4.t9 vss 15.765299f
C521 3rd_3_OTA_0.vd4.t4 vss 0.047335f
C522 3rd_3_OTA_0.vd4.t6 vss 0.414091f
C523 3rd_3_OTA_0.vd4.t5 vss 0.460228f
C524 3rd_3_OTA_0.vd4.n1 vss 2.41751f
C525 3rd_3_OTA_0.vd4.t0 vss 0.087062f
C526 3rd_3_OTA_0.vd4.t7 vss 0.087062f
C527 3rd_3_OTA_0.vd4.n2 vss 0.241817f
C528 3rd_3_OTA_0.vd4.n3 vss 1.40386f
C529 3rd_3_OTA_0.vd4.n4 vss 1.3906f
C530 3rd_3_OTA_0.vd4.t2 vss 0.042702f
C531 3rd_3_OTA_0.vd4.t3 vss 0.008706f
C532 3rd_3_OTA_0.vd4.t1 vss 0.008706f
C533 3rd_3_OTA_0.vd4.n5 vss 0.0515f
C534 a_n1236_n9479.n0 vss 0.297823f
C535 a_n1236_n9479.n1 vss 0.297439f
C536 a_n1236_n9479.n2 vss 0.29823f
C537 a_n1236_n9479.n3 vss 0.29615f
C538 a_n1236_n9479.n4 vss 0.295296f
C539 a_n1236_n9479.n5 vss 0.585351f
C540 a_n1236_n9479.n6 vss 0.294838f
C541 a_n1236_n9479.n7 vss 0.126637f
C542 a_n1236_n9479.n8 vss 0.297117f
C543 a_n1236_n9479.n9 vss 0.755844f
C544 a_n1236_n9479.n10 vss 0.293675f
C545 a_n1236_n9479.n11 vss 0.295194f
C546 a_n1236_n9479.n12 vss 0.292701f
C547 a_n1236_n9479.n13 vss 0.232375f
C548 a_n1236_n9479.t46 vss 0.036678f
C549 a_n1236_n9479.n14 vss 0.160547f
C550 a_n1236_n9479.n15 vss 0.15275f
C551 a_n1236_n9479.t6 vss 0.428407f
C552 a_n1236_n9479.n16 vss 0.188243f
C553 a_n1236_n9479.t37 vss 0.036678f
C554 a_n1236_n9479.t17 vss 0.036678f
C555 a_n1236_n9479.n17 vss 0.078298f
C556 a_n1236_n9479.n18 vss 0.188647f
C557 a_n1236_n9479.t16 vss 0.428407f
C558 a_n1236_n9479.n19 vss 0.126601f
C559 a_n1236_n9479.t30 vss 0.428407f
C560 a_n1236_n9479.n20 vss 0.191708f
C561 a_n1236_n9479.n21 vss 0.191714f
C562 a_n1236_n9479.n22 vss 0.126636f
C563 a_n1236_n9479.n23 vss 0.252394f
C564 a_n1236_n9479.n24 vss 0.235053f
C565 a_n1236_n9479.t14 vss 0.429053f
C566 a_n1236_n9479.n25 vss 0.501918f
C567 a_n1236_n9479.t15 vss 0.036678f
C568 a_n1236_n9479.t36 vss 0.036678f
C569 a_n1236_n9479.n26 vss 0.078351f
C570 a_n1236_n9479.t39 vss 0.036678f
C571 a_n1236_n9479.t3 vss 0.036678f
C572 a_n1236_n9479.n27 vss 0.078351f
C573 a_n1236_n9479.n28 vss 0.209863f
C574 a_n1236_n9479.n29 vss 0.152512f
C575 a_n1236_n9479.n30 vss 0.210635f
C576 a_n1236_n9479.t2 vss 0.428407f
C577 a_n1236_n9479.n31 vss 0.244957f
C578 a_n1236_n9479.t28 vss 0.428407f
C579 a_n1236_n9479.n32 vss 0.198133f
C580 a_n1236_n9479.n33 vss 0.152497f
C581 a_n1236_n9479.t29 vss 0.036678f
C582 a_n1236_n9479.t45 vss 0.036678f
C583 a_n1236_n9479.n34 vss 0.078351f
C584 a_n1236_n9479.t40 vss 0.036678f
C585 a_n1236_n9479.t7 vss 0.036678f
C586 a_n1236_n9479.n35 vss 0.078353f
C587 a_n1236_n9479.n36 vss 0.224428f
C588 a_n1236_n9479.n37 vss 0.194658f
C589 a_n1236_n9479.t4 vss 0.428407f
C590 a_n1236_n9479.t0 vss 0.429046f
C591 a_n1236_n9479.t21 vss 0.036678f
C592 a_n1236_n9479.t38 vss 0.036678f
C593 a_n1236_n9479.n38 vss 0.078351f
C594 a_n1236_n9479.t42 vss 0.036678f
C595 a_n1236_n9479.t1 vss 0.036678f
C596 a_n1236_n9479.n39 vss 0.078351f
C597 a_n1236_n9479.n40 vss 0.281102f
C598 a_n1236_n9479.n41 vss 0.512311f
C599 a_n1236_n9479.n42 vss 0.190453f
C600 a_n1236_n9479.t23 vss 0.036678f
C601 a_n1236_n9479.t47 vss 0.036678f
C602 a_n1236_n9479.n43 vss 0.078298f
C603 a_n1236_n9479.t34 vss 0.036678f
C604 a_n1236_n9479.t11 vss 0.036678f
C605 a_n1236_n9479.n44 vss 0.078298f
C606 a_n1236_n9479.n45 vss 0.192954f
C607 a_n1236_n9479.t24 vss 0.428407f
C608 a_n1236_n9479.n46 vss 0.126637f
C609 a_n1236_n9479.n47 vss 0.229843f
C610 a_n1236_n9479.t10 vss 0.428407f
C611 a_n1236_n9479.n48 vss 0.19241f
C612 a_n1236_n9479.n49 vss 0.196776f
C613 a_n1236_n9479.n50 vss 0.133795f
C614 a_n1236_n9479.t25 vss 0.036678f
C615 a_n1236_n9479.t32 vss 0.036678f
C616 a_n1236_n9479.n51 vss 0.078298f
C617 a_n1236_n9479.t43 vss 0.036678f
C618 a_n1236_n9479.t9 vss 0.036678f
C619 a_n1236_n9479.n52 vss 0.078298f
C620 a_n1236_n9479.t27 vss 0.036678f
C621 a_n1236_n9479.t33 vss 0.036678f
C622 a_n1236_n9479.n53 vss 0.078508f
C623 a_n1236_n9479.n54 vss 0.109851f
C624 a_n1236_n9479.n55 vss 0.128037f
C625 a_n1236_n9479.t26 vss 0.428407f
C626 a_n1236_n9479.n56 vss 0.194392f
C627 a_n1236_n9479.n57 vss 0.192707f
C628 a_n1236_n9479.t8 vss 0.428407f
C629 a_n1236_n9479.n58 vss 0.252273f
C630 a_n1236_n9479.n59 vss 0.285147f
C631 a_n1236_n9479.n60 vss 0.138692f
C632 a_n1236_n9479.n61 vss 0.126601f
C633 a_n1236_n9479.n62 vss 0.195682f
C634 a_n1236_n9479.t20 vss 0.428407f
C635 a_n1236_n9479.n63 vss 0.185109f
C636 a_n1236_n9479.n64 vss 0.213178f
C637 a_n1236_n9479.n65 vss 0.126622f
C638 a_n1236_n9479.n66 vss 0.074228f
C639 a_n1236_n9479.t41 vss 0.036678f
C640 a_n1236_n9479.t5 vss 0.036678f
C641 a_n1236_n9479.n67 vss 0.078351f
C642 a_n1236_n9479.n68 vss 0.224594f
C643 a_n1236_n9479.t19 vss 0.036678f
C644 a_n1236_n9479.t44 vss 0.036678f
C645 a_n1236_n9479.n69 vss 0.078351f
C646 a_n1236_n9479.n70 vss 0.191262f
C647 a_n1236_n9479.t18 vss 0.428407f
C648 a_n1236_n9479.n71 vss 0.181786f
C649 a_n1236_n9479.n72 vss 0.116531f
C650 a_n1236_n9479.n73 vss 0.075366f
C651 a_n1236_n9479.n74 vss 0.116443f
C652 a_n1236_n9479.n75 vss 0.160573f
C653 a_n1236_n9479.n76 vss 0.15275f
C654 a_n1236_n9479.n77 vss 0.230436f
C655 a_n1236_n9479.n78 vss 0.126601f
C656 a_n1236_n9479.n79 vss 0.188243f
C657 a_n1236_n9479.t22 vss 0.428407f
C658 a_n1236_n9479.n80 vss 0.192694f
C659 a_n1236_n9479.t12 vss 0.428407f
C660 a_n1236_n9479.n81 vss 0.191841f
C661 a_n1236_n9479.n82 vss 0.126638f
C662 a_n1236_n9479.t35 vss 0.036678f
C663 a_n1236_n9479.t13 vss 0.036678f
C664 a_n1236_n9479.n83 vss 0.078298f
C665 a_n1236_n9479.n84 vss 0.078298f
C666 a_n1236_n9479.t31 vss 0.036678f
C667 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 vss 7.77106f
C668 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 vss 5.32305f
C669 OTA_vref_0.OTA_vref_stage2_0.vref0.t32 vss 0.077096f
C670 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 vss 0.07938f
C671 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 vss 0.07938f
C672 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 vss 0.278065f
C673 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 vss 0.07938f
C674 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 vss 0.07938f
C675 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 vss 0.254416f
C676 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 vss 0.07938f
C677 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 vss 0.07938f
C678 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 vss 0.254416f
C679 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 vss 0.07938f
C680 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 vss 0.07938f
C681 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 vss 0.254416f
C682 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 vss 0.07938f
C683 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 vss 0.07938f
C684 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 vss 0.254416f
C685 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 vss 0.07938f
C686 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 vss 0.07938f
C687 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 vss 0.254416f
C688 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 vss 0.07938f
C689 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 vss 0.07938f
C690 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 vss 0.254416f
C691 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 vss 0.07938f
C692 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 vss 0.07938f
C693 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 vss 0.254416f
C694 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 vss 0.07938f
C695 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 vss 0.07938f
C696 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 vss 0.254284f
C697 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 vss 0.07938f
C698 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 vss 0.07938f
C699 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 vss 0.254416f
C700 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 vss 0.07938f
C701 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 vss 0.07938f
C702 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 vss 0.264281f
C703 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 vss 0.07938f
C704 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 vss 0.07938f
C705 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 vss 0.254416f
C706 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 vss 0.07938f
C707 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 vss 0.07938f
C708 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 vss 0.254416f
C709 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 vss 0.07938f
C710 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 vss 0.07938f
C711 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 vss 0.254416f
C712 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 vss 0.07938f
C713 OTA_vref_0.OTA_vref_stage2_0.vref0.t0 vss 0.07938f
C714 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 vss 0.254416f
C715 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 vss 0.07938f
C716 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 vss 0.07938f
C717 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 vss 0.254416f
C718 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 vss 0.072231f
C719 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 vss 0.110183f
C720 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 vss 0.109159f
C721 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 vss -3.70902f
C722 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 vss 3.98388f
C723 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 vss 0.478981f
C724 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 vss 0.480213f
C725 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 vss 1.17119f
C726 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 vss 0.305431f
C727 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 vss 0.478028f
C728 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 vss 0.234187f
C729 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 vss 0.470573f
C730 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 vss 0.478028f
C731 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 vss 0.470573f
C732 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 vss 0.478028f
C733 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 vss 0.470129f
C734 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 vss 0.478028f
C735 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 vss 0.119324f
C736 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 vss 0.391163f
C737 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 vss 0.207747f
C738 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 vss 0.305316f
C739 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 vss 0.478809f
C740 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 vss 0.222027f
C741 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 vss 0.474153f
C742 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 vss 0.478028f
C743 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 vss 0.474153f
C744 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 vss 0.478028f
C745 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 vss 0.472108f
C746 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 vss 0.478028f
C747 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 vss 0.114607f
C748 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 vss 0.358056f
C749 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 vss 0.1713f
C750 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 vss 0.305164f
C751 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 vss 0.478028f
C752 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 vss 0.234725f
C753 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 vss 0.471116f
C754 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 vss 0.478028f
C755 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 vss 0.471116f
C756 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 vss 0.478028f
C757 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 vss 0.471016f
C758 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 vss 0.478028f
C759 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 vss 0.116651f
C760 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 vss 0.391917f
C761 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 vss 0.175402f
C762 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 vss 0.305187f
C763 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 vss 0.478881f
C764 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 vss 0.232796f
C765 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 vss 0.470031f
C766 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 vss 0.478028f
C767 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 vss 0.470031f
C768 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 vss 0.478028f
C769 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 vss 0.470335f
C770 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 vss 0.478028f
C771 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 vss 0.118954f
C772 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 vss 0.357235f
C773 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 vss 0.171379f
C774 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 vss 0.305728f
C775 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 vss 0.478028f
C776 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 vss 0.231521f
C777 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 vss 0.470851f
C778 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 vss 0.478028f
C779 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 vss 0.470852f
C780 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 vss 0.478028f
C781 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 vss 0.466741f
C782 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 vss 0.478028f
C783 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 vss 0.124091f
C784 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 vss 0.391922f
C785 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 vss 0.175402f
C786 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 vss 0.478028f
C787 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 vss 0.28265f
C788 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 vss 0.46793f
C789 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 vss 0.478028f
C790 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 vss 0.240285f
C791 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 vss 0.478028f
C792 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 vss 0.46793f
C793 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 vss 0.304748f
C794 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 vss 0.478028f
C795 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 vss 0.303889f
C796 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 vss 0.157732f
C797 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 vss 0.205161f
C798 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 vss 0.171854f
C799 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 vss 0.305508f
C800 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 vss 0.478028f
C801 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 vss 0.22844f
C802 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 vss 0.473853f
C803 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 vss 0.478028f
C804 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 vss 0.473853f
C805 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 vss 0.478028f
C806 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 vss 0.473079f
C807 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 vss 0.478028f
C808 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 vss 0.113695f
C809 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 vss 0.395354f
C810 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 vss 0.17643f
C811 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 vss 0.480413f
C812 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 vss 0.478986f
C813 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 vss 1.18519f
C814 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 vss 0.383039f
C815 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 vss 0.473185f
C816 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 vss 0.215214f
C817 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 vss 0.201225f
C818 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 vss 0.215214f
C819 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 vss 0.215214f
C820 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 vss 0.184059f
C821 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 vss 0.04125f
C822 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 vss 0.041255f
C823 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 vss 1.0568f
C824 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 vss 0.444711f
C825 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 vss 0.122425f
C826 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 vss 0.110183f
C827 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 vss 0.10796f
C828 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 vss 0.122425f
C829 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 vss 0.490623f
C830 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n92 vss 0.201231f
C831 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n94 vss 0.381488f
C832 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n95 vss 0.147422f
C833 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n96 vss 0.329195f
C834 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n97 vss 0.122425f
C835 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n98 vss 0.21592f
C836 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n99 vss 0.21592f
C837 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n100 vss 0.101613f
C838 a_7434_495.n0 vss 0.6008f
C839 a_7434_495.n1 vss 0.948802f
C840 a_7434_495.n2 vss 1.1133f
C841 a_7434_495.n3 vss 0.22981f
C842 a_7434_495.n4 vss 2.01666f
C843 a_7434_495.n5 vss 0.043049f
C844 a_7434_495.n6 vss 0.034133f
C845 a_7434_495.n7 vss 2.02362f
C846 a_7434_495.n8 vss 1.9823f
C847 a_7434_495.t0 vss 0.1247f
C848 a_7434_495.t12 vss 0.105673f
C849 a_7434_495.t7 vss 0.067294f
C850 a_7434_495.t6 vss 1.20911f
C851 a_7434_495.t5 vss 0.018244f
C852 a_7434_495.t9 vss 0.018244f
C853 a_7434_495.n9 vss 0.037169f
C854 a_7434_495.n10 vss 0.069191f
C855 a_7434_495.n11 vss 0.235173f
C856 a_7434_495.t8 vss 1.21226f
C857 a_7434_495.t4 vss 1.20913f
C858 a_7434_495.t10 vss 1.20913f
C859 a_7434_495.n12 vss 1.96965f
C860 a_7434_495.t11 vss 0.067212f
C861 a_7434_495.n13 vss 0.327769f
C862 a_7434_495.n14 vss 1.14135f
C863 a_7434_495.t1 vss 0.021893f
C864 a_7434_495.t2 vss 0.021893f
C865 a_7434_495.n15 vss 0.069059f
C866 a_7434_495.n16 vss 1.00528f
C867 a_7434_495.n17 vss 1.25188f
C868 a_7434_495.t3 vss 0.116219f
C869 3rd_3_OTA_0.vd3.n0 vss 1.01087f
C870 3rd_3_OTA_0.vd3.n1 vss 1.90811f
C871 3rd_3_OTA_0.vd3.n2 vss 1.76973f
C872 3rd_3_OTA_0.vd3.n3 vss 0.035523f
C873 3rd_3_OTA_0.vd3.n4 vss 1.7787f
C874 3rd_3_OTA_0.vd3.n5 vss 1.94522f
C875 3rd_3_OTA_0.vd3.t19 vss 0.276606f
C876 3rd_3_OTA_0.vd3.t18 vss 0.276453f
C877 3rd_3_OTA_0.vd3.t13 vss 0.276526f
C878 3rd_3_OTA_0.vd3.t12 vss 0.274737f
C879 3rd_3_OTA_0.vd3.t10 vss 0.04613f
C880 3rd_3_OTA_0.vd3.t9 vss 0.04613f
C881 3rd_3_OTA_0.vd3.n6 vss 0.145431f
C882 3rd_3_OTA_0.vd3.t11 vss 0.210471f
C883 3rd_3_OTA_0.vd3.t0 vss 0.232664f
C884 3rd_3_OTA_0.vd3.n7 vss 0.615792f
C885 3rd_3_OTA_0.vd3.t4 vss 0.016281f
C886 3rd_3_OTA_0.vd3.t8 vss 0.016281f
C887 3rd_3_OTA_0.vd3.t7 vss 0.641539f
C888 3rd_3_OTA_0.vd3.t16 vss 0.641537f
C889 3rd_3_OTA_0.vd3.n8 vss 0.239118f
C890 3rd_3_OTA_0.vd3.t15 vss 0.641539f
C891 3rd_3_OTA_0.vd3.t5 vss 0.641537f
C892 3rd_3_OTA_0.vd3.n9 vss 0.239118f
C893 3rd_3_OTA_0.vd3.t6 vss 0.004613f
C894 3rd_3_OTA_0.vd3.t2 vss 0.004613f
C895 3rd_3_OTA_0.vd3.n10 vss 0.009758f
C896 3rd_3_OTA_0.vd3.t17 vss 0.641539f
C897 3rd_3_OTA_0.vd3.t1 vss 0.641537f
C898 3rd_3_OTA_0.vd3.n11 vss 0.239118f
C899 3rd_3_OTA_0.vd3.t3 vss 0.641539f
C900 3rd_3_OTA_0.vd3.t14 vss 0.641537f
C901 3rd_3_OTA_0.vd3.n12 vss 0.239118f
C902 3rd_3_OTA_0.vd3.n13 vss 1.71789f
.ends

