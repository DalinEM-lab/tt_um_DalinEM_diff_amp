magic
tech sky130A
magscale 1 2
timestamp 1741292250
<< metal1 >>
rect 26488 9458 26498 9459
rect 25886 9358 26498 9458
rect 26488 9298 26498 9358
rect 26678 9298 26688 9459
<< via1 >>
rect 26498 9298 26678 9459
<< metal2 >>
rect 11712 31140 11935 33016
rect 10935 31121 11665 31131
rect 10935 30951 11665 30961
rect 29707 24249 29886 24259
rect 27759 24069 29707 24249
rect 29707 24058 29886 24068
rect 9129 23600 9383 23610
rect 9383 23382 11835 23600
rect 11870 23594 19325 23604
rect 9129 23372 9383 23382
rect 11870 23381 19325 23391
rect 11526 21341 11683 21351
rect 11683 20968 12120 21341
rect 11526 20958 11683 20968
rect 30362 20775 30542 20785
rect 30362 17647 30542 20632
rect 30358 17477 30367 17647
rect 30537 17477 30546 17647
rect 30362 17472 30542 17477
rect 30362 13028 30542 13038
rect 13963 12273 14168 12283
rect 7845 11892 13963 12273
rect 1903 10420 2303 10430
rect 2303 10020 2701 10420
rect 7845 10381 8226 11892
rect 13963 11882 14168 11892
rect 25902 11404 26136 11414
rect 25902 10994 26136 11004
rect 7847 10380 8226 10381
rect 1903 10010 2303 10020
rect 26498 9459 26678 9469
rect 26498 9288 26678 9298
rect 30362 8230 30542 12891
rect 30362 8077 30542 8087
rect 11501 6554 11886 6563
rect 11501 5732 11886 6169
rect 11501 5347 17832 5732
rect 17447 5332 17727 5347
rect 7178 2767 7358 3098
rect 7178 2648 7358 2658
<< via2 >>
rect 10935 30961 11665 31121
rect 29707 24068 29886 24249
rect 9129 23382 9383 23600
rect 11870 23391 19325 23594
rect 11526 20968 11683 21341
rect 30362 20632 30542 20775
rect 30367 17477 30537 17647
rect 30362 12891 30542 13028
rect 13963 11892 14168 12273
rect 1903 10020 2303 10420
rect 25902 11004 26136 11404
rect 26498 9303 26678 9458
rect 30362 8087 30542 8230
rect 11501 6169 11886 6554
rect 7178 2658 7358 2767
<< metal3 >>
rect 10925 31121 11675 31126
rect 10925 30961 10935 31121
rect 11665 30961 11675 31121
rect 10925 30956 11675 30961
rect 4927 12970 5107 24434
rect 7385 13785 7565 24542
rect 29697 24249 29896 24254
rect 29697 24068 29707 24249
rect 29886 24068 29896 24249
rect 29697 24063 29896 24068
rect 9119 23600 9393 23605
rect 9119 23382 9129 23600
rect 9383 23382 9393 23600
rect 11860 23594 19335 23599
rect 11860 23391 11870 23594
rect 19325 23391 19335 23594
rect 11860 23386 19335 23391
rect 9119 23377 9393 23382
rect 11516 21341 11693 21346
rect 11516 20968 11526 21341
rect 11683 20968 11693 21341
rect 11516 20963 11693 20968
rect 30352 20775 30552 20780
rect 30352 20632 30362 20775
rect 30542 20632 30552 20775
rect 30352 20627 30552 20632
rect 30363 17652 30541 17657
rect 30362 17651 30542 17652
rect 30362 17473 30363 17651
rect 30541 17473 30542 17651
rect 30362 17472 30542 17473
rect 30363 17467 30541 17472
rect 7385 13605 11623 13785
rect 11772 13605 11782 13785
rect 30352 13028 30552 13033
rect 4927 12790 9240 12970
rect 9417 12790 9427 12970
rect 30352 12891 30362 13028
rect 30542 12891 30552 13028
rect 30352 12886 30552 12891
rect 13953 12273 14178 12278
rect 13953 11892 13963 12273
rect 14168 11892 14178 12273
rect 13953 11887 14178 11892
rect 4867 11174 4873 11559
rect 5258 11174 11886 11559
rect 1893 10420 2313 10425
rect 1893 10020 1903 10420
rect 2303 10020 2313 10420
rect 1893 10015 2313 10020
rect 11501 6559 11886 11174
rect 25892 11404 26146 11409
rect 25892 11004 25902 11404
rect 26136 11004 26146 11404
rect 25892 10999 26146 11004
rect 26488 9458 26688 9463
rect 26488 9303 26498 9458
rect 26678 9303 26688 9458
rect 26488 9298 26688 9303
rect 30352 8230 30552 8235
rect 30352 8087 30362 8230
rect 30542 8087 30552 8230
rect 30352 8082 30552 8087
rect 11496 6554 11891 6559
rect 11496 6169 11501 6554
rect 11886 6169 11891 6554
rect 11496 6164 11891 6169
rect 18663 3571 18843 5309
rect 14906 3391 18843 3571
rect 7168 2767 7368 2772
rect 7168 2658 7178 2767
rect 7358 2658 7368 2767
rect 7168 2653 7368 2658
rect 14906 1818 15086 3391
rect 19436 2805 19616 5283
rect 21894 4301 22074 5281
rect 21884 4121 21894 4301
rect 22074 4121 22084 4301
rect 21894 4119 22074 4121
rect 19426 2625 19436 2805
rect 19616 2625 19626 2805
rect 14896 1638 14906 1818
rect 15086 1638 15096 1818
<< via3 >>
rect 10935 30961 11665 31121
rect 29707 24068 29886 24249
rect 9129 23382 9383 23600
rect 11870 23391 19325 23594
rect 11526 20968 11683 21341
rect 30362 20632 30542 20775
rect 30363 17647 30541 17651
rect 30363 17477 30367 17647
rect 30367 17477 30537 17647
rect 30537 17477 30541 17647
rect 30363 17473 30541 17477
rect 11623 13605 11772 13785
rect 9240 12790 9417 12970
rect 30362 12891 30542 13028
rect 13963 11892 14168 12273
rect 4873 11174 5258 11559
rect 1903 10020 2303 10420
rect 25902 11004 26136 11404
rect 26498 9303 26678 9458
rect 30362 8087 30542 8230
rect 7178 2658 7358 2767
rect 21894 4121 22074 4301
rect 19436 2625 19616 2805
rect 14906 1638 15086 1818
<< metal4 >>
rect 400 43919 800 44152
rect 400 43282 2000 43919
rect 400 25519 800 43282
rect 31400 33199 31800 44152
rect 11470 31122 11930 33197
rect 14344 32876 31800 33199
rect 14500 32798 31800 32876
rect 14502 32797 31800 32798
rect 10934 31121 11930 31122
rect 10934 30961 10935 31121
rect 11665 30961 11930 31121
rect 10934 30960 11930 30961
rect 11470 30794 11930 30960
rect 31400 30560 31800 32797
rect 31399 30160 31800 30560
rect 31400 28175 31800 30160
rect 29046 27621 31800 28175
rect 400 25327 3015 25519
rect 400 25119 2980 25327
rect 400 23600 800 25119
rect 29706 24249 29887 24250
rect 29706 24068 29707 24249
rect 29886 24069 30542 24249
rect 29886 24068 29887 24069
rect 29706 24067 29887 24068
rect 9128 23600 9384 23601
rect 400 23382 9129 23600
rect 9383 23382 9384 23600
rect 19288 23595 20764 23600
rect 11869 23594 20764 23595
rect 11869 23391 11870 23594
rect 19325 23391 20764 23594
rect 11869 23390 20764 23391
rect 19288 23384 20764 23390
rect 400 11559 800 23382
rect 8157 21341 8530 23382
rect 9128 23381 9384 23382
rect 11525 21341 11684 21342
rect 8157 20968 11526 21341
rect 11683 20968 11684 21341
rect 11525 20967 11684 20968
rect 30362 20776 30542 24069
rect 30361 20775 30543 20776
rect 30361 20632 30362 20775
rect 30542 20632 30543 20775
rect 30361 20631 30543 20632
rect 31400 19852 31800 27621
rect 31401 19365 31800 19852
rect 31400 19044 31800 19365
rect 29076 18490 31800 19044
rect 30362 17651 30542 17652
rect 30362 17473 30363 17651
rect 30541 17473 30542 17651
rect 11622 13785 11773 13786
rect 11622 13605 11623 13785
rect 11772 13605 13005 13785
rect 11622 13604 11773 13605
rect 9239 12970 9418 12971
rect 9239 12790 9240 12970
rect 9417 12790 10547 12970
rect 9239 12789 9418 12790
rect 4872 11559 5259 11560
rect 400 11174 4873 11559
rect 5258 11174 5259 11559
rect 400 10420 800 11174
rect 4872 11173 5259 11174
rect 1902 10420 2304 10421
rect 400 10020 1903 10420
rect 2303 10020 2304 10420
rect 400 1000 800 10020
rect 1902 10019 2304 10020
rect 10367 2805 10547 12790
rect 12825 4301 13005 13605
rect 30362 13029 30542 17473
rect 30361 13028 30543 13029
rect 30361 12891 30362 13028
rect 30542 12891 30543 13028
rect 30361 12890 30543 12891
rect 13962 12273 14169 12274
rect 13962 11892 13963 12273
rect 14168 11892 27933 12273
rect 13962 11891 14169 11892
rect 25901 11404 26137 11405
rect 27552 11404 27933 11892
rect 31400 11404 31800 18490
rect 25901 11004 25902 11404
rect 26136 11004 31800 11404
rect 25901 11003 26137 11004
rect 26497 9458 26679 9459
rect 26497 9303 26498 9458
rect 26678 9303 26679 9458
rect 26497 9302 26679 9303
rect 21893 4301 22075 4302
rect 12825 4121 21894 4301
rect 22074 4121 22814 4301
rect 21893 4120 22075 4121
rect 19435 2805 19617 2806
rect 7177 2767 7359 2768
rect 7177 2658 7178 2767
rect 7358 2658 7359 2767
rect 7177 2657 7359 2658
rect 7178 1683 7358 2657
rect 10367 2625 19436 2805
rect 19616 2625 19617 2805
rect 14905 1818 15087 1819
rect 7178 1503 11222 1683
rect 14905 1638 14906 1818
rect 15086 1638 15087 1818
rect 14905 1637 15087 1638
rect 11042 338 11222 1503
rect 11041 199 11222 338
rect 11042 0 11222 199
rect 14906 0 15086 1637
rect 18770 0 18950 2625
rect 19435 2624 19617 2625
rect 22634 0 22814 4121
rect 26498 0 26678 9302
rect 30361 8230 30543 8231
rect 30361 8087 30362 8230
rect 30542 8087 30543 8230
rect 30361 8086 30543 8087
rect 30362 0 30542 8086
rect 31400 1000 31800 11004
use 3_OTA  3_OTA_0 ~/Project_tinytape/magic/mag/3_OTA
timestamp 1741224942
transform 1 0 13614 0 1 25385
box -10693 -10528 15660 7813
use BGR_BJT_vref  BGR_BJT_vref_0 ~/Project_tinytape/magic/mag/OTA_vref
timestamp 1740770860
transform 0 -1 8258 -1 0 10672
box 0 0 7872 5648
use Diff_amp  Diff_amp_0 ~/Project_tinytape/magic/mag/OTA_stage1
timestamp 1740708554
transform 1 0 9041 0 1 31945
box 0 0 1 1
use diff_final_v0  diff_final_v0_0 ~/Project_tinytape/magic/mag/OTA_stage1
timestamp 1738105933
transform 1 0 6731 0 1 8024
box 10993 -2832 19171 3381
<< labels >>
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 31401 1000 31800 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 1000 800 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
