magic
tech sky130A
magscale 1 2
timestamp 1738270755
<< error_p >>
rect -244 -200 244 200
<< nwell >>
rect -244 -200 244 200
<< pmoslvt >>
rect -150 -100 150 100
<< pdiff >>
rect -208 88 -150 100
rect -208 -88 -196 88
rect -162 -88 -150 88
rect -208 -100 -150 -88
rect 150 88 208 100
rect 150 -88 162 88
rect 196 -88 208 88
rect 150 -100 208 -88
<< pdiffc >>
rect -196 -88 -162 88
rect 162 -88 196 88
<< poly >>
rect -150 181 150 197
rect -150 147 -134 181
rect 134 147 150 181
rect -150 100 150 147
rect -150 -147 150 -100
rect -150 -181 -134 -147
rect 134 -181 150 -147
rect -150 -197 150 -181
<< polycont >>
rect -134 147 134 181
rect -134 -181 134 -147
<< locali >>
rect -150 147 -134 181
rect 134 147 150 181
rect -196 88 -162 104
rect -196 -104 -162 -88
rect 162 88 196 104
rect 162 -104 196 -88
rect -150 -181 -134 -147
rect 134 -181 150 -147
<< viali >>
rect -134 147 134 181
rect -196 -88 -162 88
rect 162 -88 196 88
rect -134 -181 134 -147
<< metal1 >>
rect -146 181 146 187
rect -146 147 -134 181
rect 134 147 146 181
rect -146 141 146 147
rect -202 88 -156 100
rect -202 -88 -196 88
rect -162 -88 -156 88
rect -202 -100 -156 -88
rect 156 88 202 100
rect 156 -88 162 88
rect 196 -88 202 88
rect 156 -100 202 -88
rect -146 -147 146 -141
rect -146 -181 -134 -147
rect 134 -181 146 -147
rect -146 -187 146 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 1.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
