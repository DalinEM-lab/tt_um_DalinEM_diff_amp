magic
tech sky130A
magscale 1 2
timestamp 1739140642
<< nwell >>
rect 13 998 1197 999
rect 13 367 2028 998
rect 2371 368 3163 1006
rect 3661 368 4453 1006
rect 4951 368 5743 1006
rect 17 366 2028 367
rect 6247 355 7620 990
<< pwell >>
rect -1 4363 6841 5607
rect -1 4359 2159 4363
rect 2191 4359 6841 4363
rect -1 4313 6841 4359
rect -1 4310 2157 4313
rect 2190 4310 6841 4313
rect -1 2493 6841 4310
rect 53 2294 1393 2447
rect 53 1260 206 2294
rect 1240 1260 1393 2294
rect 53 1107 1393 1260
rect 1960 1051 7634 1898
<< nbase >>
rect 206 1260 1240 2294
<< pmoslvt >>
rect 247 686 647 786
rect 705 686 1105 786
rect 1372 586 1572 786
rect 1630 586 1830 786
rect 2567 587 2967 787
rect 3857 587 4257 787
rect 5147 587 5547 787
rect 6437 587 6837 787
rect 7018 587 7418 787
<< nmoslvt >>
rect 365 4391 565 5191
rect 623 4391 823 5191
rect 881 4391 1081 5191
rect 1139 4391 1339 5191
rect 1397 4391 1597 5191
rect 1655 4391 1855 5191
rect 1913 4391 2113 5191
rect 2171 4391 2371 5191
rect 2429 4391 2629 5191
rect 2687 4391 2887 5191
rect 2945 4391 3145 5191
rect 3203 4391 3403 5191
rect 3461 4391 3661 5191
rect 3719 4391 3919 5191
rect 3977 4391 4177 5191
rect 4235 4391 4435 5191
rect 4493 4391 4693 5191
rect 4751 4391 4951 5191
rect 5009 4391 5209 5191
rect 5267 4391 5467 5191
rect 5525 4391 5725 5191
rect 5783 4391 5983 5191
rect 6041 4391 6241 5191
rect 6299 4391 6499 5191
rect 365 2910 565 3710
rect 623 2910 823 3710
rect 881 2910 1081 3710
rect 1139 2910 1339 3710
rect 1397 2910 1597 3710
rect 1655 2910 1855 3710
rect 1913 2910 2113 3710
rect 2171 2910 2371 3710
rect 2429 2910 2629 3710
rect 2687 2910 2887 3710
rect 2945 2910 3145 3710
rect 3203 2910 3403 3710
rect 3461 2910 3661 3710
rect 3719 2910 3919 3710
rect 3977 2910 4177 3710
rect 4235 2910 4435 3710
rect 4493 2910 4693 3710
rect 4751 2910 4951 3710
rect 5009 2910 5209 3710
rect 5267 2910 5467 3710
rect 5525 2910 5725 3710
rect 5783 2910 5983 3710
rect 6041 2910 6241 3710
rect 6299 2910 6499 3710
rect 2251 1374 2451 1574
rect 2509 1374 2709 1574
rect 2767 1374 2967 1574
rect 3025 1374 3225 1574
rect 3283 1374 3483 1574
rect 3541 1374 3741 1574
rect 3799 1374 3999 1574
rect 4057 1374 4257 1574
rect 4315 1374 4515 1574
rect 4573 1374 4773 1574
rect 4831 1374 5031 1574
rect 5089 1374 5289 1574
rect 5347 1374 5547 1574
rect 5605 1374 5805 1574
rect 5863 1374 6063 1574
rect 6121 1374 6321 1574
rect 6379 1374 6579 1574
rect 6637 1374 6837 1574
rect 6895 1374 7095 1574
rect 7153 1374 7353 1574
<< ndiff >>
rect 307 5179 365 5191
rect 307 4403 319 5179
rect 353 4403 365 5179
rect 307 4391 365 4403
rect 565 5179 623 5191
rect 565 4403 577 5179
rect 611 4403 623 5179
rect 565 4391 623 4403
rect 823 5179 881 5191
rect 823 4403 835 5179
rect 869 4403 881 5179
rect 823 4391 881 4403
rect 1081 5179 1139 5191
rect 1081 4403 1093 5179
rect 1127 4403 1139 5179
rect 1081 4391 1139 4403
rect 1339 5179 1397 5191
rect 1339 4403 1351 5179
rect 1385 4403 1397 5179
rect 1339 4391 1397 4403
rect 1597 5179 1655 5191
rect 1597 4403 1609 5179
rect 1643 4403 1655 5179
rect 1597 4391 1655 4403
rect 1855 5179 1913 5191
rect 1855 4403 1867 5179
rect 1901 4403 1913 5179
rect 1855 4391 1913 4403
rect 2113 5179 2171 5191
rect 2113 4403 2125 5179
rect 2159 4403 2171 5179
rect 2113 4391 2171 4403
rect 2371 5179 2429 5191
rect 2371 4403 2383 5179
rect 2417 4403 2429 5179
rect 2371 4391 2429 4403
rect 2629 5179 2687 5191
rect 2629 4403 2641 5179
rect 2675 4403 2687 5179
rect 2629 4391 2687 4403
rect 2887 5179 2945 5191
rect 2887 4403 2899 5179
rect 2933 4403 2945 5179
rect 2887 4391 2945 4403
rect 3145 5179 3203 5191
rect 3145 4403 3157 5179
rect 3191 4403 3203 5179
rect 3145 4391 3203 4403
rect 3403 5179 3461 5191
rect 3403 4403 3415 5179
rect 3449 4403 3461 5179
rect 3403 4391 3461 4403
rect 3661 5179 3719 5191
rect 3661 4403 3673 5179
rect 3707 4403 3719 5179
rect 3661 4391 3719 4403
rect 3919 5179 3977 5191
rect 3919 4403 3931 5179
rect 3965 4403 3977 5179
rect 3919 4391 3977 4403
rect 4177 5179 4235 5191
rect 4177 4403 4189 5179
rect 4223 4403 4235 5179
rect 4177 4391 4235 4403
rect 4435 5179 4493 5191
rect 4435 4403 4447 5179
rect 4481 4403 4493 5179
rect 4435 4391 4493 4403
rect 4693 5179 4751 5191
rect 4693 4403 4705 5179
rect 4739 4403 4751 5179
rect 4693 4391 4751 4403
rect 4951 5179 5009 5191
rect 4951 4403 4963 5179
rect 4997 4403 5009 5179
rect 4951 4391 5009 4403
rect 5209 5179 5267 5191
rect 5209 4403 5221 5179
rect 5255 4403 5267 5179
rect 5209 4391 5267 4403
rect 5467 5179 5525 5191
rect 5467 4403 5479 5179
rect 5513 4403 5525 5179
rect 5467 4391 5525 4403
rect 5725 5179 5783 5191
rect 5725 4403 5737 5179
rect 5771 4403 5783 5179
rect 5725 4391 5783 4403
rect 5983 5179 6041 5191
rect 5983 4403 5995 5179
rect 6029 4403 6041 5179
rect 5983 4391 6041 4403
rect 6241 5179 6299 5191
rect 6241 4403 6253 5179
rect 6287 4403 6299 5179
rect 6241 4391 6299 4403
rect 6499 5179 6557 5191
rect 6499 4403 6511 5179
rect 6545 4403 6557 5179
rect 6499 4391 6557 4403
rect 307 3698 365 3710
rect 307 2922 319 3698
rect 353 2922 365 3698
rect 307 2910 365 2922
rect 565 3698 623 3710
rect 565 2922 577 3698
rect 611 2922 623 3698
rect 565 2910 623 2922
rect 823 3698 881 3710
rect 823 2922 835 3698
rect 869 2922 881 3698
rect 823 2910 881 2922
rect 1081 3698 1139 3710
rect 1081 2922 1093 3698
rect 1127 2922 1139 3698
rect 1081 2910 1139 2922
rect 1339 3698 1397 3710
rect 1339 2922 1351 3698
rect 1385 2922 1397 3698
rect 1339 2910 1397 2922
rect 1597 3698 1655 3710
rect 1597 2922 1609 3698
rect 1643 2922 1655 3698
rect 1597 2910 1655 2922
rect 1855 3698 1913 3710
rect 1855 2922 1867 3698
rect 1901 2922 1913 3698
rect 1855 2910 1913 2922
rect 2113 3698 2171 3710
rect 2113 2922 2125 3698
rect 2159 2922 2171 3698
rect 2113 2910 2171 2922
rect 2371 3698 2429 3710
rect 2371 2922 2383 3698
rect 2417 2922 2429 3698
rect 2371 2910 2429 2922
rect 2629 3698 2687 3710
rect 2629 2922 2641 3698
rect 2675 2922 2687 3698
rect 2629 2910 2687 2922
rect 2887 3698 2945 3710
rect 2887 2922 2899 3698
rect 2933 2922 2945 3698
rect 2887 2910 2945 2922
rect 3145 3698 3203 3710
rect 3145 2922 3157 3698
rect 3191 2922 3203 3698
rect 3145 2910 3203 2922
rect 3403 3698 3461 3710
rect 3403 2922 3415 3698
rect 3449 2922 3461 3698
rect 3403 2910 3461 2922
rect 3661 3698 3719 3710
rect 3661 2922 3673 3698
rect 3707 2922 3719 3698
rect 3661 2910 3719 2922
rect 3919 3698 3977 3710
rect 3919 2922 3931 3698
rect 3965 2922 3977 3698
rect 3919 2910 3977 2922
rect 4177 3698 4235 3710
rect 4177 2922 4189 3698
rect 4223 2922 4235 3698
rect 4177 2910 4235 2922
rect 4435 3698 4493 3710
rect 4435 2922 4447 3698
rect 4481 2922 4493 3698
rect 4435 2910 4493 2922
rect 4693 3698 4751 3710
rect 4693 2922 4705 3698
rect 4739 2922 4751 3698
rect 4693 2910 4751 2922
rect 4951 3698 5009 3710
rect 4951 2922 4963 3698
rect 4997 2922 5009 3698
rect 4951 2910 5009 2922
rect 5209 3698 5267 3710
rect 5209 2922 5221 3698
rect 5255 2922 5267 3698
rect 5209 2910 5267 2922
rect 5467 3698 5525 3710
rect 5467 2922 5479 3698
rect 5513 2922 5525 3698
rect 5467 2910 5525 2922
rect 5725 3698 5783 3710
rect 5725 2922 5737 3698
rect 5771 2922 5783 3698
rect 5725 2910 5783 2922
rect 5983 3698 6041 3710
rect 5983 2922 5995 3698
rect 6029 2922 6041 3698
rect 5983 2910 6041 2922
rect 6241 3698 6299 3710
rect 6241 2922 6253 3698
rect 6287 2922 6299 3698
rect 6241 2910 6299 2922
rect 6499 3698 6557 3710
rect 6499 2922 6511 3698
rect 6545 2922 6557 3698
rect 6499 2910 6557 2922
rect 2193 1562 2251 1574
rect 2193 1386 2205 1562
rect 2239 1386 2251 1562
rect 2193 1374 2251 1386
rect 2451 1562 2509 1574
rect 2451 1386 2463 1562
rect 2497 1386 2509 1562
rect 2451 1374 2509 1386
rect 2709 1562 2767 1574
rect 2709 1386 2721 1562
rect 2755 1386 2767 1562
rect 2709 1374 2767 1386
rect 2967 1562 3025 1574
rect 2967 1386 2979 1562
rect 3013 1386 3025 1562
rect 2967 1374 3025 1386
rect 3225 1562 3283 1574
rect 3225 1386 3237 1562
rect 3271 1386 3283 1562
rect 3225 1374 3283 1386
rect 3483 1562 3541 1574
rect 3483 1386 3495 1562
rect 3529 1386 3541 1562
rect 3483 1374 3541 1386
rect 3741 1562 3799 1574
rect 3741 1386 3753 1562
rect 3787 1386 3799 1562
rect 3741 1374 3799 1386
rect 3999 1562 4057 1574
rect 3999 1386 4011 1562
rect 4045 1386 4057 1562
rect 3999 1374 4057 1386
rect 4257 1562 4315 1574
rect 4257 1386 4269 1562
rect 4303 1386 4315 1562
rect 4257 1374 4315 1386
rect 4515 1562 4573 1574
rect 4515 1386 4527 1562
rect 4561 1386 4573 1562
rect 4515 1374 4573 1386
rect 4773 1562 4831 1574
rect 4773 1386 4785 1562
rect 4819 1386 4831 1562
rect 4773 1374 4831 1386
rect 5031 1562 5089 1574
rect 5031 1386 5043 1562
rect 5077 1386 5089 1562
rect 5031 1374 5089 1386
rect 5289 1562 5347 1574
rect 5289 1386 5301 1562
rect 5335 1386 5347 1562
rect 5289 1374 5347 1386
rect 5547 1562 5605 1574
rect 5547 1386 5559 1562
rect 5593 1386 5605 1562
rect 5547 1374 5605 1386
rect 5805 1562 5863 1574
rect 5805 1386 5817 1562
rect 5851 1386 5863 1562
rect 5805 1374 5863 1386
rect 6063 1562 6121 1574
rect 6063 1386 6075 1562
rect 6109 1386 6121 1562
rect 6063 1374 6121 1386
rect 6321 1562 6379 1574
rect 6321 1386 6333 1562
rect 6367 1386 6379 1562
rect 6321 1374 6379 1386
rect 6579 1562 6637 1574
rect 6579 1386 6591 1562
rect 6625 1386 6637 1562
rect 6579 1374 6637 1386
rect 6837 1562 6895 1574
rect 6837 1386 6849 1562
rect 6883 1386 6895 1562
rect 6837 1374 6895 1386
rect 7095 1562 7153 1574
rect 7095 1386 7107 1562
rect 7141 1386 7153 1562
rect 7095 1374 7153 1386
rect 7353 1562 7411 1574
rect 7353 1386 7365 1562
rect 7399 1386 7411 1562
rect 7353 1374 7411 1386
<< pdiff >>
rect 383 2065 1063 2117
rect 383 2031 437 2065
rect 471 2031 527 2065
rect 561 2031 617 2065
rect 651 2031 707 2065
rect 741 2031 797 2065
rect 831 2031 887 2065
rect 921 2031 977 2065
rect 1011 2031 1063 2065
rect 383 1975 1063 2031
rect 383 1941 437 1975
rect 471 1941 527 1975
rect 561 1941 617 1975
rect 651 1941 707 1975
rect 741 1941 797 1975
rect 831 1941 887 1975
rect 921 1941 977 1975
rect 1011 1941 1063 1975
rect 383 1885 1063 1941
rect 383 1851 437 1885
rect 471 1851 527 1885
rect 561 1851 617 1885
rect 651 1851 707 1885
rect 741 1851 797 1885
rect 831 1851 887 1885
rect 921 1851 977 1885
rect 1011 1851 1063 1885
rect 383 1795 1063 1851
rect 383 1761 437 1795
rect 471 1761 527 1795
rect 561 1761 617 1795
rect 651 1761 707 1795
rect 741 1761 797 1795
rect 831 1761 887 1795
rect 921 1761 977 1795
rect 1011 1761 1063 1795
rect 383 1705 1063 1761
rect 383 1671 437 1705
rect 471 1671 527 1705
rect 561 1671 617 1705
rect 651 1671 707 1705
rect 741 1671 797 1705
rect 831 1671 887 1705
rect 921 1671 977 1705
rect 1011 1671 1063 1705
rect 383 1615 1063 1671
rect 383 1581 437 1615
rect 471 1581 527 1615
rect 561 1581 617 1615
rect 651 1581 707 1615
rect 741 1581 797 1615
rect 831 1581 887 1615
rect 921 1581 977 1615
rect 1011 1581 1063 1615
rect 383 1525 1063 1581
rect 383 1491 437 1525
rect 471 1491 527 1525
rect 561 1491 617 1525
rect 651 1491 707 1525
rect 741 1491 797 1525
rect 831 1491 887 1525
rect 921 1491 977 1525
rect 1011 1491 1063 1525
rect 383 1437 1063 1491
rect 189 774 247 786
rect 189 698 201 774
rect 235 698 247 774
rect 189 686 247 698
rect 647 774 705 786
rect 647 698 659 774
rect 693 698 705 774
rect 647 686 705 698
rect 1105 774 1163 786
rect 1105 698 1117 774
rect 1151 698 1163 774
rect 1105 686 1163 698
rect 1314 774 1372 786
rect 1314 598 1326 774
rect 1360 598 1372 774
rect 1314 586 1372 598
rect 1572 774 1630 786
rect 1572 598 1584 774
rect 1618 598 1630 774
rect 1572 586 1630 598
rect 1830 774 1888 786
rect 1830 598 1842 774
rect 1876 598 1888 774
rect 1830 586 1888 598
rect 2509 775 2567 787
rect 2509 599 2521 775
rect 2555 599 2567 775
rect 2509 587 2567 599
rect 2967 775 3025 787
rect 2967 599 2979 775
rect 3013 599 3025 775
rect 2967 587 3025 599
rect 3799 775 3857 787
rect 3799 599 3811 775
rect 3845 599 3857 775
rect 3799 587 3857 599
rect 4257 775 4315 787
rect 4257 599 4269 775
rect 4303 599 4315 775
rect 4257 587 4315 599
rect 5089 775 5147 787
rect 5089 599 5101 775
rect 5135 599 5147 775
rect 5089 587 5147 599
rect 5547 775 5605 787
rect 5547 599 5559 775
rect 5593 599 5605 775
rect 5547 587 5605 599
rect 6379 775 6437 787
rect 6379 599 6391 775
rect 6425 599 6437 775
rect 6379 587 6437 599
rect 6837 775 6895 787
rect 6837 599 6849 775
rect 6883 599 6895 775
rect 6837 587 6895 599
rect 6960 775 7018 787
rect 6960 599 6972 775
rect 7006 599 7018 775
rect 6960 587 7018 599
rect 7418 775 7476 787
rect 7418 599 7430 775
rect 7464 599 7476 775
rect 7418 587 7476 599
<< ndiffc >>
rect 319 4403 353 5179
rect 577 4403 611 5179
rect 835 4403 869 5179
rect 1093 4403 1127 5179
rect 1351 4403 1385 5179
rect 1609 4403 1643 5179
rect 1867 4403 1901 5179
rect 2125 4403 2159 5179
rect 2383 4403 2417 5179
rect 2641 4403 2675 5179
rect 2899 4403 2933 5179
rect 3157 4403 3191 5179
rect 3415 4403 3449 5179
rect 3673 4403 3707 5179
rect 3931 4403 3965 5179
rect 4189 4403 4223 5179
rect 4447 4403 4481 5179
rect 4705 4403 4739 5179
rect 4963 4403 4997 5179
rect 5221 4403 5255 5179
rect 5479 4403 5513 5179
rect 5737 4403 5771 5179
rect 5995 4403 6029 5179
rect 6253 4403 6287 5179
rect 6511 4403 6545 5179
rect 319 2922 353 3698
rect 577 2922 611 3698
rect 835 2922 869 3698
rect 1093 2922 1127 3698
rect 1351 2922 1385 3698
rect 1609 2922 1643 3698
rect 1867 2922 1901 3698
rect 2125 2922 2159 3698
rect 2383 2922 2417 3698
rect 2641 2922 2675 3698
rect 2899 2922 2933 3698
rect 3157 2922 3191 3698
rect 3415 2922 3449 3698
rect 3673 2922 3707 3698
rect 3931 2922 3965 3698
rect 4189 2922 4223 3698
rect 4447 2922 4481 3698
rect 4705 2922 4739 3698
rect 4963 2922 4997 3698
rect 5221 2922 5255 3698
rect 5479 2922 5513 3698
rect 5737 2922 5771 3698
rect 5995 2922 6029 3698
rect 6253 2922 6287 3698
rect 6511 2922 6545 3698
rect 2205 1386 2239 1562
rect 2463 1386 2497 1562
rect 2721 1386 2755 1562
rect 2979 1386 3013 1562
rect 3237 1386 3271 1562
rect 3495 1386 3529 1562
rect 3753 1386 3787 1562
rect 4011 1386 4045 1562
rect 4269 1386 4303 1562
rect 4527 1386 4561 1562
rect 4785 1386 4819 1562
rect 5043 1386 5077 1562
rect 5301 1386 5335 1562
rect 5559 1386 5593 1562
rect 5817 1386 5851 1562
rect 6075 1386 6109 1562
rect 6333 1386 6367 1562
rect 6591 1386 6625 1562
rect 6849 1386 6883 1562
rect 7107 1386 7141 1562
rect 7365 1386 7399 1562
<< pdiffc >>
rect 437 2031 471 2065
rect 527 2031 561 2065
rect 617 2031 651 2065
rect 707 2031 741 2065
rect 797 2031 831 2065
rect 887 2031 921 2065
rect 977 2031 1011 2065
rect 437 1941 471 1975
rect 527 1941 561 1975
rect 617 1941 651 1975
rect 707 1941 741 1975
rect 797 1941 831 1975
rect 887 1941 921 1975
rect 977 1941 1011 1975
rect 437 1851 471 1885
rect 527 1851 561 1885
rect 617 1851 651 1885
rect 707 1851 741 1885
rect 797 1851 831 1885
rect 887 1851 921 1885
rect 977 1851 1011 1885
rect 437 1761 471 1795
rect 527 1761 561 1795
rect 617 1761 651 1795
rect 707 1761 741 1795
rect 797 1761 831 1795
rect 887 1761 921 1795
rect 977 1761 1011 1795
rect 437 1671 471 1705
rect 527 1671 561 1705
rect 617 1671 651 1705
rect 707 1671 741 1705
rect 797 1671 831 1705
rect 887 1671 921 1705
rect 977 1671 1011 1705
rect 437 1581 471 1615
rect 527 1581 561 1615
rect 617 1581 651 1615
rect 707 1581 741 1615
rect 797 1581 831 1615
rect 887 1581 921 1615
rect 977 1581 1011 1615
rect 437 1491 471 1525
rect 527 1491 561 1525
rect 617 1491 651 1525
rect 707 1491 741 1525
rect 797 1491 831 1525
rect 887 1491 921 1525
rect 977 1491 1011 1525
rect 201 698 235 774
rect 659 698 693 774
rect 1117 698 1151 774
rect 1326 598 1360 774
rect 1584 598 1618 774
rect 1842 598 1876 774
rect 2521 599 2555 775
rect 2979 599 3013 775
rect 3811 599 3845 775
rect 4269 599 4303 775
rect 5101 599 5135 775
rect 5559 599 5593 775
rect 6391 599 6425 775
rect 6849 599 6883 775
rect 6972 599 7006 775
rect 7430 599 7464 775
<< psubdiff >>
rect 113 5433 173 5467
rect 6629 5433 6689 5467
rect 113 5407 147 5433
rect 6655 5407 6689 5433
rect 113 2672 147 2698
rect 6655 2672 6689 2698
rect 113 2638 173 2672
rect 6629 2638 6689 2672
rect 79 2386 1367 2421
rect 79 2363 209 2386
rect 79 2329 113 2363
rect 147 2352 209 2363
rect 243 2352 299 2386
rect 333 2352 389 2386
rect 423 2352 479 2386
rect 513 2352 569 2386
rect 603 2352 659 2386
rect 693 2352 749 2386
rect 783 2352 839 2386
rect 873 2352 929 2386
rect 963 2352 1019 2386
rect 1053 2352 1109 2386
rect 1143 2352 1199 2386
rect 1233 2363 1367 2386
rect 1233 2352 1300 2363
rect 147 2329 1300 2352
rect 1334 2329 1367 2363
rect 79 2320 1367 2329
rect 79 2273 180 2320
rect 79 2239 113 2273
rect 147 2239 180 2273
rect 1266 2273 1367 2320
rect 79 2183 180 2239
rect 79 2149 113 2183
rect 147 2149 180 2183
rect 79 2093 180 2149
rect 79 2059 113 2093
rect 147 2059 180 2093
rect 79 2003 180 2059
rect 79 1969 113 2003
rect 147 1969 180 2003
rect 79 1913 180 1969
rect 79 1879 113 1913
rect 147 1879 180 1913
rect 79 1823 180 1879
rect 79 1789 113 1823
rect 147 1789 180 1823
rect 79 1733 180 1789
rect 79 1699 113 1733
rect 147 1699 180 1733
rect 79 1643 180 1699
rect 79 1609 113 1643
rect 147 1609 180 1643
rect 79 1553 180 1609
rect 79 1519 113 1553
rect 147 1519 180 1553
rect 79 1463 180 1519
rect 79 1429 113 1463
rect 147 1429 180 1463
rect 79 1373 180 1429
rect 79 1339 113 1373
rect 147 1339 180 1373
rect 79 1283 180 1339
rect 1266 2239 1300 2273
rect 1334 2239 1367 2273
rect 1266 2183 1367 2239
rect 1266 2149 1300 2183
rect 1334 2149 1367 2183
rect 1266 2093 1367 2149
rect 1266 2059 1300 2093
rect 1334 2059 1367 2093
rect 1266 2003 1367 2059
rect 1266 1969 1300 2003
rect 1334 1969 1367 2003
rect 1266 1913 1367 1969
rect 1266 1879 1300 1913
rect 1334 1879 1367 1913
rect 1266 1823 1367 1879
rect 1266 1789 1300 1823
rect 1334 1789 1367 1823
rect 1266 1733 1367 1789
rect 1266 1699 1300 1733
rect 1334 1699 1367 1733
rect 1266 1643 1367 1699
rect 1266 1609 1300 1643
rect 1334 1609 1367 1643
rect 1266 1553 1367 1609
rect 1266 1519 1300 1553
rect 1334 1519 1367 1553
rect 1266 1463 1367 1519
rect 1266 1429 1300 1463
rect 1334 1429 1367 1463
rect 1266 1373 1367 1429
rect 1266 1339 1300 1373
rect 1334 1339 1367 1373
rect 79 1249 113 1283
rect 147 1249 180 1283
rect 79 1234 180 1249
rect 1266 1283 1367 1339
rect 1266 1249 1300 1283
rect 1334 1249 1367 1283
rect 1266 1234 1367 1249
rect 79 1199 1367 1234
rect 79 1165 209 1199
rect 243 1165 299 1199
rect 333 1165 389 1199
rect 423 1165 479 1199
rect 513 1165 569 1199
rect 603 1165 659 1199
rect 693 1165 749 1199
rect 783 1165 839 1199
rect 873 1165 929 1199
rect 963 1165 1019 1199
rect 1053 1165 1109 1199
rect 1143 1165 1199 1199
rect 1233 1165 1367 1199
rect 79 1133 1367 1165
rect 2038 1786 2098 1820
rect 7506 1786 7566 1820
rect 2038 1760 2072 1786
rect 7532 1760 7566 1786
rect 2038 1152 2072 1178
rect 7532 1152 7566 1178
rect 2038 1118 2098 1152
rect 7506 1118 7566 1152
<< nsubdiff >>
rect 242 2239 1204 2258
rect 242 2205 373 2239
rect 407 2205 463 2239
rect 497 2205 553 2239
rect 587 2205 643 2239
rect 677 2205 733 2239
rect 767 2205 823 2239
rect 857 2205 913 2239
rect 947 2205 1003 2239
rect 1037 2205 1093 2239
rect 1127 2205 1204 2239
rect 242 2186 1204 2205
rect 242 2182 314 2186
rect 242 2148 261 2182
rect 295 2148 314 2182
rect 242 2092 314 2148
rect 1132 2163 1204 2186
rect 1132 2129 1151 2163
rect 1185 2129 1204 2163
rect 242 2058 261 2092
rect 295 2058 314 2092
rect 242 2002 314 2058
rect 242 1968 261 2002
rect 295 1968 314 2002
rect 242 1912 314 1968
rect 242 1878 261 1912
rect 295 1878 314 1912
rect 242 1822 314 1878
rect 242 1788 261 1822
rect 295 1788 314 1822
rect 242 1732 314 1788
rect 242 1698 261 1732
rect 295 1698 314 1732
rect 242 1642 314 1698
rect 242 1608 261 1642
rect 295 1608 314 1642
rect 242 1552 314 1608
rect 242 1518 261 1552
rect 295 1518 314 1552
rect 242 1462 314 1518
rect 242 1428 261 1462
rect 295 1428 314 1462
rect 1132 2073 1204 2129
rect 1132 2039 1151 2073
rect 1185 2039 1204 2073
rect 1132 1983 1204 2039
rect 1132 1949 1151 1983
rect 1185 1949 1204 1983
rect 1132 1893 1204 1949
rect 1132 1859 1151 1893
rect 1185 1859 1204 1893
rect 1132 1803 1204 1859
rect 1132 1769 1151 1803
rect 1185 1769 1204 1803
rect 1132 1713 1204 1769
rect 1132 1679 1151 1713
rect 1185 1679 1204 1713
rect 1132 1623 1204 1679
rect 1132 1589 1151 1623
rect 1185 1589 1204 1623
rect 1132 1533 1204 1589
rect 1132 1499 1151 1533
rect 1185 1499 1204 1533
rect 1132 1443 1204 1499
rect 242 1368 314 1428
rect 1132 1409 1151 1443
rect 1185 1409 1204 1443
rect 1132 1368 1204 1409
rect 242 1349 1204 1368
rect 242 1315 339 1349
rect 373 1315 429 1349
rect 463 1315 519 1349
rect 553 1315 609 1349
rect 643 1315 699 1349
rect 733 1315 789 1349
rect 823 1315 879 1349
rect 913 1315 969 1349
rect 1003 1315 1059 1349
rect 1093 1315 1204 1349
rect 242 1296 1204 1315
rect 51 912 239 960
rect 1347 912 1604 960
rect 1881 912 1992 960
rect 51 793 103 912
rect 1943 877 1992 912
rect 51 462 103 557
rect 1943 462 1992 498
rect 51 410 199 462
rect 1874 410 1992 462
rect 2407 936 2503 970
rect 3031 936 3127 970
rect 2407 874 2441 936
rect 3093 874 3127 936
rect 2407 438 2441 500
rect 3093 438 3127 500
rect 2407 404 2503 438
rect 3031 404 3127 438
rect 3697 936 3793 970
rect 4321 936 4417 970
rect 3697 874 3731 936
rect 4383 874 4417 936
rect 3697 438 3731 500
rect 4383 438 4417 500
rect 3697 404 3793 438
rect 4321 404 4417 438
rect 4987 936 5083 970
rect 5611 936 5707 970
rect 4987 874 5021 936
rect 5673 874 5707 936
rect 4987 438 5021 500
rect 5673 438 5707 500
rect 4987 404 5083 438
rect 5611 404 5707 438
rect 6290 912 6350 946
rect 7514 912 7574 946
rect 6290 886 6324 912
rect 7540 886 7574 912
rect 6290 436 6324 462
rect 7540 436 7574 462
rect 6290 402 6350 436
rect 7514 402 7574 436
<< psubdiffcont >>
rect 173 5433 6629 5467
rect 113 2698 147 5407
rect 6655 2698 6689 5407
rect 173 2638 6629 2672
rect 113 2329 147 2363
rect 209 2352 243 2386
rect 299 2352 333 2386
rect 389 2352 423 2386
rect 479 2352 513 2386
rect 569 2352 603 2386
rect 659 2352 693 2386
rect 749 2352 783 2386
rect 839 2352 873 2386
rect 929 2352 963 2386
rect 1019 2352 1053 2386
rect 1109 2352 1143 2386
rect 1199 2352 1233 2386
rect 1300 2329 1334 2363
rect 113 2239 147 2273
rect 113 2149 147 2183
rect 113 2059 147 2093
rect 113 1969 147 2003
rect 113 1879 147 1913
rect 113 1789 147 1823
rect 113 1699 147 1733
rect 113 1609 147 1643
rect 113 1519 147 1553
rect 113 1429 147 1463
rect 113 1339 147 1373
rect 1300 2239 1334 2273
rect 1300 2149 1334 2183
rect 1300 2059 1334 2093
rect 1300 1969 1334 2003
rect 1300 1879 1334 1913
rect 1300 1789 1334 1823
rect 1300 1699 1334 1733
rect 1300 1609 1334 1643
rect 1300 1519 1334 1553
rect 1300 1429 1334 1463
rect 1300 1339 1334 1373
rect 113 1249 147 1283
rect 1300 1249 1334 1283
rect 209 1165 243 1199
rect 299 1165 333 1199
rect 389 1165 423 1199
rect 479 1165 513 1199
rect 569 1165 603 1199
rect 659 1165 693 1199
rect 749 1165 783 1199
rect 839 1165 873 1199
rect 929 1165 963 1199
rect 1019 1165 1053 1199
rect 1109 1165 1143 1199
rect 1199 1165 1233 1199
rect 2098 1786 7506 1820
rect 2038 1178 2072 1760
rect 7532 1178 7566 1760
rect 2098 1118 7506 1152
<< nsubdiffcont >>
rect 373 2205 407 2239
rect 463 2205 497 2239
rect 553 2205 587 2239
rect 643 2205 677 2239
rect 733 2205 767 2239
rect 823 2205 857 2239
rect 913 2205 947 2239
rect 1003 2205 1037 2239
rect 1093 2205 1127 2239
rect 261 2148 295 2182
rect 1151 2129 1185 2163
rect 261 2058 295 2092
rect 261 1968 295 2002
rect 261 1878 295 1912
rect 261 1788 295 1822
rect 261 1698 295 1732
rect 261 1608 295 1642
rect 261 1518 295 1552
rect 261 1428 295 1462
rect 1151 2039 1185 2073
rect 1151 1949 1185 1983
rect 1151 1859 1185 1893
rect 1151 1769 1185 1803
rect 1151 1679 1185 1713
rect 1151 1589 1185 1623
rect 1151 1499 1185 1533
rect 1151 1409 1185 1443
rect 339 1315 373 1349
rect 429 1315 463 1349
rect 519 1315 553 1349
rect 609 1315 643 1349
rect 699 1315 733 1349
rect 789 1315 823 1349
rect 879 1315 913 1349
rect 969 1315 1003 1349
rect 1059 1315 1093 1349
rect 239 912 1347 960
rect 1604 912 1881 960
rect 51 557 103 793
rect 1943 498 1992 877
rect 199 410 1874 462
rect 2503 936 3031 970
rect 2407 500 2441 874
rect 3093 500 3127 874
rect 2503 404 3031 438
rect 3793 936 4321 970
rect 3697 500 3731 874
rect 4383 500 4417 874
rect 3793 404 4321 438
rect 5083 936 5611 970
rect 4987 500 5021 874
rect 5673 500 5707 874
rect 5083 404 5611 438
rect 6350 912 7514 946
rect 6290 462 6324 886
rect 7540 462 7574 886
rect 6350 402 7514 436
<< poly >>
rect 365 5263 565 5279
rect 365 5229 381 5263
rect 549 5229 565 5263
rect 365 5191 565 5229
rect 623 5263 823 5279
rect 623 5229 639 5263
rect 807 5229 823 5263
rect 623 5191 823 5229
rect 881 5263 1081 5279
rect 881 5229 897 5263
rect 1065 5229 1081 5263
rect 881 5191 1081 5229
rect 1139 5263 1339 5279
rect 1139 5229 1155 5263
rect 1323 5229 1339 5263
rect 1139 5191 1339 5229
rect 1397 5263 1597 5279
rect 1397 5229 1413 5263
rect 1581 5229 1597 5263
rect 1397 5191 1597 5229
rect 1655 5263 1855 5279
rect 1655 5229 1671 5263
rect 1839 5229 1855 5263
rect 1655 5191 1855 5229
rect 1913 5263 2113 5279
rect 1913 5229 1929 5263
rect 2097 5229 2113 5263
rect 1913 5191 2113 5229
rect 2171 5263 2371 5279
rect 2171 5229 2187 5263
rect 2355 5229 2371 5263
rect 2171 5191 2371 5229
rect 2429 5263 2629 5279
rect 2429 5229 2445 5263
rect 2613 5229 2629 5263
rect 2429 5191 2629 5229
rect 2687 5263 2887 5279
rect 2687 5229 2703 5263
rect 2871 5229 2887 5263
rect 2687 5191 2887 5229
rect 2945 5263 3145 5279
rect 2945 5229 2961 5263
rect 3129 5229 3145 5263
rect 2945 5191 3145 5229
rect 3203 5263 3403 5279
rect 3203 5229 3219 5263
rect 3387 5229 3403 5263
rect 3203 5191 3403 5229
rect 3461 5263 3661 5279
rect 3461 5229 3477 5263
rect 3645 5229 3661 5263
rect 3461 5191 3661 5229
rect 3719 5263 3919 5279
rect 3719 5229 3735 5263
rect 3903 5229 3919 5263
rect 3719 5191 3919 5229
rect 3977 5263 4177 5279
rect 3977 5229 3993 5263
rect 4161 5229 4177 5263
rect 3977 5191 4177 5229
rect 4235 5263 4435 5279
rect 4235 5229 4251 5263
rect 4419 5229 4435 5263
rect 4235 5191 4435 5229
rect 4493 5263 4693 5279
rect 4493 5229 4509 5263
rect 4677 5229 4693 5263
rect 4493 5191 4693 5229
rect 4751 5263 4951 5279
rect 4751 5229 4767 5263
rect 4935 5229 4951 5263
rect 4751 5191 4951 5229
rect 5009 5263 5209 5279
rect 5009 5229 5025 5263
rect 5193 5229 5209 5263
rect 5009 5191 5209 5229
rect 5267 5263 5467 5279
rect 5267 5229 5283 5263
rect 5451 5229 5467 5263
rect 5267 5191 5467 5229
rect 5525 5263 5725 5279
rect 5525 5229 5541 5263
rect 5709 5229 5725 5263
rect 5525 5191 5725 5229
rect 5783 5263 5983 5279
rect 5783 5229 5799 5263
rect 5967 5229 5983 5263
rect 5783 5191 5983 5229
rect 6041 5263 6241 5279
rect 6041 5229 6057 5263
rect 6225 5229 6241 5263
rect 6041 5191 6241 5229
rect 6299 5263 6499 5279
rect 6299 5229 6315 5263
rect 6483 5229 6499 5263
rect 6299 5191 6499 5229
rect 365 4353 565 4391
rect 365 4319 381 4353
rect 549 4319 565 4353
rect 365 4303 565 4319
rect 623 4353 823 4391
rect 623 4319 639 4353
rect 807 4319 823 4353
rect 623 4303 823 4319
rect 881 4353 1081 4391
rect 881 4319 897 4353
rect 1065 4319 1081 4353
rect 881 4303 1081 4319
rect 1139 4353 1339 4391
rect 1139 4319 1155 4353
rect 1323 4319 1339 4353
rect 1139 4303 1339 4319
rect 1397 4353 1597 4391
rect 1397 4319 1413 4353
rect 1581 4319 1597 4353
rect 1397 4303 1597 4319
rect 1655 4353 1855 4391
rect 1655 4319 1671 4353
rect 1839 4319 1855 4353
rect 1655 4303 1855 4319
rect 1913 4353 2113 4391
rect 1913 4319 1929 4353
rect 2097 4319 2113 4353
rect 1913 4303 2113 4319
rect 2171 4353 2371 4391
rect 2171 4319 2187 4353
rect 2355 4319 2371 4353
rect 2171 4303 2371 4319
rect 2429 4353 2629 4391
rect 2429 4319 2445 4353
rect 2613 4319 2629 4353
rect 2429 4303 2629 4319
rect 2687 4353 2887 4391
rect 2687 4319 2703 4353
rect 2871 4319 2887 4353
rect 2687 4303 2887 4319
rect 2945 4353 3145 4391
rect 2945 4319 2961 4353
rect 3129 4319 3145 4353
rect 2945 4303 3145 4319
rect 3203 4353 3403 4391
rect 3203 4319 3219 4353
rect 3387 4319 3403 4353
rect 3203 4303 3403 4319
rect 3461 4353 3661 4391
rect 3461 4319 3477 4353
rect 3645 4319 3661 4353
rect 3461 4303 3661 4319
rect 3719 4353 3919 4391
rect 3719 4319 3735 4353
rect 3903 4319 3919 4353
rect 3719 4303 3919 4319
rect 3977 4353 4177 4391
rect 3977 4319 3993 4353
rect 4161 4319 4177 4353
rect 3977 4303 4177 4319
rect 4235 4353 4435 4391
rect 4235 4319 4251 4353
rect 4419 4319 4435 4353
rect 4235 4303 4435 4319
rect 4493 4353 4693 4391
rect 4493 4319 4509 4353
rect 4677 4319 4693 4353
rect 4493 4303 4693 4319
rect 4751 4353 4951 4391
rect 4751 4319 4767 4353
rect 4935 4319 4951 4353
rect 4751 4303 4951 4319
rect 5009 4353 5209 4391
rect 5009 4319 5025 4353
rect 5193 4319 5209 4353
rect 5009 4303 5209 4319
rect 5267 4353 5467 4391
rect 5267 4319 5283 4353
rect 5451 4319 5467 4353
rect 5267 4303 5467 4319
rect 5525 4353 5725 4391
rect 5525 4319 5541 4353
rect 5709 4319 5725 4353
rect 5525 4303 5725 4319
rect 5783 4353 5983 4391
rect 5783 4319 5799 4353
rect 5967 4319 5983 4353
rect 5783 4303 5983 4319
rect 6041 4353 6241 4391
rect 6041 4319 6057 4353
rect 6225 4319 6241 4353
rect 6041 4303 6241 4319
rect 6299 4353 6499 4391
rect 6299 4319 6315 4353
rect 6483 4319 6499 4353
rect 6299 4303 6499 4319
rect 365 3782 565 3798
rect 365 3748 381 3782
rect 549 3748 565 3782
rect 365 3710 565 3748
rect 623 3782 823 3798
rect 623 3748 639 3782
rect 807 3748 823 3782
rect 623 3710 823 3748
rect 881 3782 1081 3798
rect 881 3748 897 3782
rect 1065 3748 1081 3782
rect 881 3710 1081 3748
rect 1139 3782 1339 3798
rect 1139 3748 1155 3782
rect 1323 3748 1339 3782
rect 1139 3710 1339 3748
rect 1397 3782 1597 3798
rect 1397 3748 1413 3782
rect 1581 3748 1597 3782
rect 1397 3710 1597 3748
rect 1655 3782 1855 3798
rect 1655 3748 1671 3782
rect 1839 3748 1855 3782
rect 1655 3710 1855 3748
rect 1913 3782 2113 3798
rect 1913 3748 1929 3782
rect 2097 3748 2113 3782
rect 1913 3710 2113 3748
rect 2171 3782 2371 3798
rect 2171 3748 2187 3782
rect 2355 3748 2371 3782
rect 2171 3710 2371 3748
rect 2429 3782 2629 3798
rect 2429 3748 2445 3782
rect 2613 3748 2629 3782
rect 2429 3710 2629 3748
rect 2687 3782 2887 3798
rect 2687 3748 2703 3782
rect 2871 3748 2887 3782
rect 2687 3710 2887 3748
rect 2945 3782 3145 3798
rect 2945 3748 2961 3782
rect 3129 3748 3145 3782
rect 2945 3710 3145 3748
rect 3203 3782 3403 3798
rect 3203 3748 3219 3782
rect 3387 3748 3403 3782
rect 3203 3710 3403 3748
rect 3461 3782 3661 3798
rect 3461 3748 3477 3782
rect 3645 3748 3661 3782
rect 3461 3710 3661 3748
rect 3719 3782 3919 3798
rect 3719 3748 3735 3782
rect 3903 3748 3919 3782
rect 3719 3710 3919 3748
rect 3977 3782 4177 3798
rect 3977 3748 3993 3782
rect 4161 3748 4177 3782
rect 3977 3710 4177 3748
rect 4235 3782 4435 3798
rect 4235 3748 4251 3782
rect 4419 3748 4435 3782
rect 4235 3710 4435 3748
rect 4493 3782 4693 3798
rect 4493 3748 4509 3782
rect 4677 3748 4693 3782
rect 4493 3710 4693 3748
rect 4751 3782 4951 3798
rect 4751 3748 4767 3782
rect 4935 3748 4951 3782
rect 4751 3710 4951 3748
rect 5009 3782 5209 3798
rect 5009 3748 5025 3782
rect 5193 3748 5209 3782
rect 5009 3710 5209 3748
rect 5267 3782 5467 3798
rect 5267 3748 5283 3782
rect 5451 3748 5467 3782
rect 5267 3710 5467 3748
rect 5525 3782 5725 3798
rect 5525 3748 5541 3782
rect 5709 3748 5725 3782
rect 5525 3710 5725 3748
rect 5783 3782 5983 3798
rect 5783 3748 5799 3782
rect 5967 3748 5983 3782
rect 5783 3710 5983 3748
rect 6041 3782 6241 3798
rect 6041 3748 6057 3782
rect 6225 3748 6241 3782
rect 6041 3710 6241 3748
rect 6299 3782 6499 3798
rect 6299 3748 6315 3782
rect 6483 3748 6499 3782
rect 6299 3710 6499 3748
rect 365 2872 565 2910
rect 365 2838 381 2872
rect 549 2838 565 2872
rect 365 2822 565 2838
rect 623 2872 823 2910
rect 623 2838 639 2872
rect 807 2838 823 2872
rect 623 2822 823 2838
rect 881 2872 1081 2910
rect 881 2838 897 2872
rect 1065 2838 1081 2872
rect 881 2822 1081 2838
rect 1139 2872 1339 2910
rect 1139 2838 1155 2872
rect 1323 2838 1339 2872
rect 1139 2822 1339 2838
rect 1397 2872 1597 2910
rect 1397 2838 1413 2872
rect 1581 2838 1597 2872
rect 1397 2822 1597 2838
rect 1655 2872 1855 2910
rect 1655 2838 1671 2872
rect 1839 2838 1855 2872
rect 1655 2822 1855 2838
rect 1913 2872 2113 2910
rect 1913 2838 1929 2872
rect 2097 2838 2113 2872
rect 1913 2822 2113 2838
rect 2171 2872 2371 2910
rect 2171 2838 2187 2872
rect 2355 2838 2371 2872
rect 2171 2822 2371 2838
rect 2429 2872 2629 2910
rect 2429 2838 2445 2872
rect 2613 2838 2629 2872
rect 2429 2822 2629 2838
rect 2687 2872 2887 2910
rect 2687 2838 2703 2872
rect 2871 2838 2887 2872
rect 2687 2822 2887 2838
rect 2945 2872 3145 2910
rect 2945 2838 2961 2872
rect 3129 2838 3145 2872
rect 2945 2822 3145 2838
rect 3203 2872 3403 2910
rect 3203 2838 3219 2872
rect 3387 2838 3403 2872
rect 3203 2822 3403 2838
rect 3461 2872 3661 2910
rect 3461 2838 3477 2872
rect 3645 2838 3661 2872
rect 3461 2822 3661 2838
rect 3719 2872 3919 2910
rect 3719 2838 3735 2872
rect 3903 2838 3919 2872
rect 3719 2822 3919 2838
rect 3977 2872 4177 2910
rect 3977 2838 3993 2872
rect 4161 2838 4177 2872
rect 3977 2822 4177 2838
rect 4235 2872 4435 2910
rect 4235 2838 4251 2872
rect 4419 2838 4435 2872
rect 4235 2822 4435 2838
rect 4493 2872 4693 2910
rect 4493 2838 4509 2872
rect 4677 2838 4693 2872
rect 4493 2822 4693 2838
rect 4751 2872 4951 2910
rect 4751 2838 4767 2872
rect 4935 2838 4951 2872
rect 4751 2822 4951 2838
rect 5009 2872 5209 2910
rect 5009 2838 5025 2872
rect 5193 2838 5209 2872
rect 5009 2822 5209 2838
rect 5267 2872 5467 2910
rect 5267 2838 5283 2872
rect 5451 2838 5467 2872
rect 5267 2822 5467 2838
rect 5525 2872 5725 2910
rect 5525 2838 5541 2872
rect 5709 2838 5725 2872
rect 5525 2822 5725 2838
rect 5783 2872 5983 2910
rect 5783 2838 5799 2872
rect 5967 2838 5983 2872
rect 5783 2822 5983 2838
rect 6041 2872 6241 2910
rect 6041 2838 6057 2872
rect 6225 2838 6241 2872
rect 6041 2822 6241 2838
rect 6299 2872 6499 2910
rect 6299 2838 6315 2872
rect 6483 2838 6499 2872
rect 6299 2822 6499 2838
rect 2251 1646 2451 1662
rect 2251 1612 2267 1646
rect 2435 1612 2451 1646
rect 2251 1574 2451 1612
rect 2509 1646 2709 1662
rect 2509 1612 2525 1646
rect 2693 1612 2709 1646
rect 2509 1574 2709 1612
rect 2767 1646 2967 1662
rect 2767 1612 2783 1646
rect 2951 1612 2967 1646
rect 2767 1574 2967 1612
rect 3025 1646 3225 1662
rect 3025 1612 3041 1646
rect 3209 1612 3225 1646
rect 3025 1574 3225 1612
rect 3283 1646 3483 1662
rect 3283 1612 3299 1646
rect 3467 1612 3483 1646
rect 3283 1574 3483 1612
rect 3541 1646 3741 1662
rect 3541 1612 3557 1646
rect 3725 1612 3741 1646
rect 3541 1574 3741 1612
rect 3799 1646 3999 1662
rect 3799 1612 3815 1646
rect 3983 1612 3999 1646
rect 3799 1574 3999 1612
rect 4057 1646 4257 1662
rect 4057 1612 4073 1646
rect 4241 1612 4257 1646
rect 4057 1574 4257 1612
rect 4315 1646 4515 1662
rect 4315 1612 4331 1646
rect 4499 1612 4515 1646
rect 4315 1574 4515 1612
rect 4573 1646 4773 1662
rect 4573 1612 4589 1646
rect 4757 1612 4773 1646
rect 4573 1574 4773 1612
rect 4831 1646 5031 1662
rect 4831 1612 4847 1646
rect 5015 1612 5031 1646
rect 4831 1574 5031 1612
rect 5089 1646 5289 1662
rect 5089 1612 5105 1646
rect 5273 1612 5289 1646
rect 5089 1574 5289 1612
rect 5347 1646 5547 1662
rect 5347 1612 5363 1646
rect 5531 1612 5547 1646
rect 5347 1574 5547 1612
rect 5605 1646 5805 1662
rect 5605 1612 5621 1646
rect 5789 1612 5805 1646
rect 5605 1574 5805 1612
rect 5863 1646 6063 1662
rect 5863 1612 5879 1646
rect 6047 1612 6063 1646
rect 5863 1574 6063 1612
rect 6121 1646 6321 1662
rect 6121 1612 6137 1646
rect 6305 1612 6321 1646
rect 6121 1574 6321 1612
rect 6379 1646 6579 1662
rect 6379 1612 6395 1646
rect 6563 1612 6579 1646
rect 6379 1574 6579 1612
rect 6637 1646 6837 1662
rect 6637 1612 6653 1646
rect 6821 1612 6837 1646
rect 6637 1574 6837 1612
rect 6895 1646 7095 1662
rect 6895 1612 6911 1646
rect 7079 1612 7095 1646
rect 6895 1574 7095 1612
rect 7153 1646 7353 1662
rect 7153 1612 7169 1646
rect 7337 1612 7353 1646
rect 7153 1574 7353 1612
rect 2251 1336 2451 1374
rect 2251 1302 2267 1336
rect 2435 1302 2451 1336
rect 2251 1286 2451 1302
rect 2509 1336 2709 1374
rect 2509 1302 2525 1336
rect 2693 1302 2709 1336
rect 2509 1286 2709 1302
rect 2767 1336 2967 1374
rect 2767 1302 2783 1336
rect 2951 1302 2967 1336
rect 2767 1286 2967 1302
rect 3025 1336 3225 1374
rect 3025 1302 3041 1336
rect 3209 1302 3225 1336
rect 3025 1286 3225 1302
rect 3283 1336 3483 1374
rect 3283 1302 3299 1336
rect 3467 1302 3483 1336
rect 3283 1286 3483 1302
rect 3541 1336 3741 1374
rect 3541 1302 3557 1336
rect 3725 1302 3741 1336
rect 3541 1286 3741 1302
rect 3799 1336 3999 1374
rect 3799 1302 3815 1336
rect 3983 1302 3999 1336
rect 3799 1286 3999 1302
rect 4057 1336 4257 1374
rect 4057 1302 4073 1336
rect 4241 1302 4257 1336
rect 4057 1286 4257 1302
rect 4315 1336 4515 1374
rect 4315 1302 4331 1336
rect 4499 1302 4515 1336
rect 4315 1286 4515 1302
rect 4573 1336 4773 1374
rect 4573 1302 4589 1336
rect 4757 1302 4773 1336
rect 4573 1286 4773 1302
rect 4831 1336 5031 1374
rect 4831 1302 4847 1336
rect 5015 1302 5031 1336
rect 4831 1286 5031 1302
rect 5089 1336 5289 1374
rect 5089 1302 5105 1336
rect 5273 1302 5289 1336
rect 5089 1286 5289 1302
rect 5347 1336 5547 1374
rect 5347 1302 5363 1336
rect 5531 1302 5547 1336
rect 5347 1286 5547 1302
rect 5605 1336 5805 1374
rect 5605 1302 5621 1336
rect 5789 1302 5805 1336
rect 5605 1286 5805 1302
rect 5863 1336 6063 1374
rect 5863 1302 5879 1336
rect 6047 1302 6063 1336
rect 5863 1286 6063 1302
rect 6121 1336 6321 1374
rect 6121 1302 6137 1336
rect 6305 1302 6321 1336
rect 6121 1286 6321 1302
rect 6379 1336 6579 1374
rect 6379 1302 6395 1336
rect 6563 1302 6579 1336
rect 6379 1286 6579 1302
rect 6637 1336 6837 1374
rect 6637 1302 6653 1336
rect 6821 1302 6837 1336
rect 6637 1286 6837 1302
rect 6895 1336 7095 1374
rect 6895 1302 6911 1336
rect 7079 1302 7095 1336
rect 6895 1286 7095 1302
rect 7153 1336 7353 1374
rect 7153 1302 7169 1336
rect 7337 1302 7353 1336
rect 7153 1286 7353 1302
rect 247 867 647 883
rect 247 833 263 867
rect 631 833 647 867
rect 247 786 647 833
rect 705 867 1105 883
rect 705 833 721 867
rect 1089 833 1105 867
rect 705 786 1105 833
rect 1372 867 1572 883
rect 1372 833 1388 867
rect 1556 833 1572 867
rect 1372 786 1572 833
rect 1630 867 1830 883
rect 1630 833 1646 867
rect 1814 833 1830 867
rect 1630 786 1830 833
rect 247 639 647 686
rect 247 605 263 639
rect 631 605 647 639
rect 247 589 647 605
rect 705 639 1105 686
rect 705 605 721 639
rect 1089 605 1105 639
rect 705 589 1105 605
rect 1372 539 1572 586
rect 1372 505 1388 539
rect 1556 505 1572 539
rect 1372 489 1572 505
rect 1630 539 1830 586
rect 1630 505 1646 539
rect 1814 505 1830 539
rect 1630 489 1830 505
rect 2567 868 2967 884
rect 2567 834 2583 868
rect 2951 834 2967 868
rect 2567 787 2967 834
rect 2567 540 2967 587
rect 2567 506 2583 540
rect 2951 506 2967 540
rect 2567 490 2967 506
rect 3857 868 4257 884
rect 3857 834 3873 868
rect 4241 834 4257 868
rect 3857 787 4257 834
rect 3857 540 4257 587
rect 3857 506 3873 540
rect 4241 506 4257 540
rect 3857 490 4257 506
rect 5147 868 5547 884
rect 5147 834 5163 868
rect 5531 834 5547 868
rect 5147 787 5547 834
rect 5147 540 5547 587
rect 5147 506 5163 540
rect 5531 506 5547 540
rect 5147 490 5547 506
rect 6437 868 6837 884
rect 6437 834 6453 868
rect 6821 834 6837 868
rect 6437 787 6837 834
rect 7018 868 7418 884
rect 7018 834 7034 868
rect 7402 834 7418 868
rect 7018 787 7418 834
rect 6437 540 6837 587
rect 6437 506 6453 540
rect 6821 506 6837 540
rect 6437 490 6837 506
rect 7018 540 7418 587
rect 7018 506 7034 540
rect 7402 506 7418 540
rect 7018 490 7418 506
<< polycont >>
rect 381 5229 549 5263
rect 639 5229 807 5263
rect 897 5229 1065 5263
rect 1155 5229 1323 5263
rect 1413 5229 1581 5263
rect 1671 5229 1839 5263
rect 1929 5229 2097 5263
rect 2187 5229 2355 5263
rect 2445 5229 2613 5263
rect 2703 5229 2871 5263
rect 2961 5229 3129 5263
rect 3219 5229 3387 5263
rect 3477 5229 3645 5263
rect 3735 5229 3903 5263
rect 3993 5229 4161 5263
rect 4251 5229 4419 5263
rect 4509 5229 4677 5263
rect 4767 5229 4935 5263
rect 5025 5229 5193 5263
rect 5283 5229 5451 5263
rect 5541 5229 5709 5263
rect 5799 5229 5967 5263
rect 6057 5229 6225 5263
rect 6315 5229 6483 5263
rect 381 4319 549 4353
rect 639 4319 807 4353
rect 897 4319 1065 4353
rect 1155 4319 1323 4353
rect 1413 4319 1581 4353
rect 1671 4319 1839 4353
rect 1929 4319 2097 4353
rect 2187 4319 2355 4353
rect 2445 4319 2613 4353
rect 2703 4319 2871 4353
rect 2961 4319 3129 4353
rect 3219 4319 3387 4353
rect 3477 4319 3645 4353
rect 3735 4319 3903 4353
rect 3993 4319 4161 4353
rect 4251 4319 4419 4353
rect 4509 4319 4677 4353
rect 4767 4319 4935 4353
rect 5025 4319 5193 4353
rect 5283 4319 5451 4353
rect 5541 4319 5709 4353
rect 5799 4319 5967 4353
rect 6057 4319 6225 4353
rect 6315 4319 6483 4353
rect 381 3748 549 3782
rect 639 3748 807 3782
rect 897 3748 1065 3782
rect 1155 3748 1323 3782
rect 1413 3748 1581 3782
rect 1671 3748 1839 3782
rect 1929 3748 2097 3782
rect 2187 3748 2355 3782
rect 2445 3748 2613 3782
rect 2703 3748 2871 3782
rect 2961 3748 3129 3782
rect 3219 3748 3387 3782
rect 3477 3748 3645 3782
rect 3735 3748 3903 3782
rect 3993 3748 4161 3782
rect 4251 3748 4419 3782
rect 4509 3748 4677 3782
rect 4767 3748 4935 3782
rect 5025 3748 5193 3782
rect 5283 3748 5451 3782
rect 5541 3748 5709 3782
rect 5799 3748 5967 3782
rect 6057 3748 6225 3782
rect 6315 3748 6483 3782
rect 381 2838 549 2872
rect 639 2838 807 2872
rect 897 2838 1065 2872
rect 1155 2838 1323 2872
rect 1413 2838 1581 2872
rect 1671 2838 1839 2872
rect 1929 2838 2097 2872
rect 2187 2838 2355 2872
rect 2445 2838 2613 2872
rect 2703 2838 2871 2872
rect 2961 2838 3129 2872
rect 3219 2838 3387 2872
rect 3477 2838 3645 2872
rect 3735 2838 3903 2872
rect 3993 2838 4161 2872
rect 4251 2838 4419 2872
rect 4509 2838 4677 2872
rect 4767 2838 4935 2872
rect 5025 2838 5193 2872
rect 5283 2838 5451 2872
rect 5541 2838 5709 2872
rect 5799 2838 5967 2872
rect 6057 2838 6225 2872
rect 6315 2838 6483 2872
rect 2267 1612 2435 1646
rect 2525 1612 2693 1646
rect 2783 1612 2951 1646
rect 3041 1612 3209 1646
rect 3299 1612 3467 1646
rect 3557 1612 3725 1646
rect 3815 1612 3983 1646
rect 4073 1612 4241 1646
rect 4331 1612 4499 1646
rect 4589 1612 4757 1646
rect 4847 1612 5015 1646
rect 5105 1612 5273 1646
rect 5363 1612 5531 1646
rect 5621 1612 5789 1646
rect 5879 1612 6047 1646
rect 6137 1612 6305 1646
rect 6395 1612 6563 1646
rect 6653 1612 6821 1646
rect 6911 1612 7079 1646
rect 7169 1612 7337 1646
rect 2267 1302 2435 1336
rect 2525 1302 2693 1336
rect 2783 1302 2951 1336
rect 3041 1302 3209 1336
rect 3299 1302 3467 1336
rect 3557 1302 3725 1336
rect 3815 1302 3983 1336
rect 4073 1302 4241 1336
rect 4331 1302 4499 1336
rect 4589 1302 4757 1336
rect 4847 1302 5015 1336
rect 5105 1302 5273 1336
rect 5363 1302 5531 1336
rect 5621 1302 5789 1336
rect 5879 1302 6047 1336
rect 6137 1302 6305 1336
rect 6395 1302 6563 1336
rect 6653 1302 6821 1336
rect 6911 1302 7079 1336
rect 7169 1302 7337 1336
rect 263 833 631 867
rect 721 833 1089 867
rect 1388 833 1556 867
rect 1646 833 1814 867
rect 263 605 631 639
rect 721 605 1089 639
rect 1388 505 1556 539
rect 1646 505 1814 539
rect 2583 834 2951 868
rect 2583 506 2951 540
rect 3873 834 4241 868
rect 3873 506 4241 540
rect 5163 834 5531 868
rect 5163 506 5531 540
rect 6453 834 6821 868
rect 7034 834 7402 868
rect 6453 506 6821 540
rect 7034 506 7402 540
<< locali >>
rect -6 5604 6712 5682
rect -6 5430 97 5604
rect 6675 5430 6712 5604
rect -6 5407 6712 5430
rect -6 5348 113 5407
rect 147 5348 6655 5407
rect -6 5321 100 5348
rect 81 5196 100 5321
rect 154 5321 6655 5348
rect 154 5196 173 5321
rect 365 5229 381 5263
rect 549 5229 565 5263
rect 623 5229 639 5263
rect 807 5229 823 5263
rect 881 5229 897 5263
rect 1065 5229 1081 5263
rect 1139 5229 1155 5263
rect 1323 5229 1339 5263
rect 1397 5229 1413 5263
rect 1581 5229 1597 5263
rect 1655 5229 1671 5263
rect 1839 5229 1855 5263
rect 1913 5229 1929 5263
rect 2097 5229 2113 5263
rect 2171 5229 2187 5263
rect 2355 5229 2371 5263
rect 2429 5229 2445 5263
rect 2613 5229 2629 5263
rect 2687 5229 2703 5263
rect 2871 5229 2887 5263
rect 2945 5229 2961 5263
rect 3129 5229 3145 5263
rect 3203 5229 3219 5263
rect 3387 5229 3403 5263
rect 3461 5229 3477 5263
rect 3645 5229 3661 5263
rect 3719 5229 3735 5263
rect 3903 5229 3919 5263
rect 3977 5229 3993 5263
rect 4161 5229 4177 5263
rect 4235 5229 4251 5263
rect 4419 5229 4435 5263
rect 4493 5229 4509 5263
rect 4677 5229 4693 5263
rect 4751 5229 4767 5263
rect 4935 5229 4951 5263
rect 5009 5229 5025 5263
rect 5193 5229 5209 5263
rect 5267 5229 5283 5263
rect 5451 5229 5467 5263
rect 5525 5229 5541 5263
rect 5709 5229 5725 5263
rect 5783 5229 5799 5263
rect 5967 5229 5983 5263
rect 6041 5229 6057 5263
rect 6225 5229 6241 5263
rect 6299 5229 6315 5263
rect 6483 5229 6499 5263
rect 81 4358 113 5196
rect 147 4358 173 5196
rect 319 5179 353 5195
rect 319 4387 353 4403
rect 577 5179 611 5195
rect 577 4387 611 4403
rect 835 5179 869 5195
rect 835 4387 869 4403
rect 1093 5179 1127 5195
rect 1093 4387 1127 4403
rect 1351 5179 1385 5195
rect 1351 4387 1385 4403
rect 1609 5179 1643 5195
rect 1609 4387 1643 4403
rect 1867 5179 1901 5195
rect 1867 4387 1901 4403
rect 2125 5179 2159 5195
rect 2125 4387 2159 4403
rect 2383 5179 2417 5195
rect 2383 4387 2417 4403
rect 2641 5179 2675 5195
rect 2641 4387 2675 4403
rect 2899 5179 2933 5195
rect 2899 4387 2933 4403
rect 3157 5179 3191 5195
rect 3157 4387 3191 4403
rect 3415 5179 3449 5195
rect 3415 4387 3449 4403
rect 3673 5179 3707 5195
rect 3673 4387 3707 4403
rect 3931 5179 3965 5195
rect 3931 4387 3965 4403
rect 4189 5179 4223 5195
rect 4189 4387 4223 4403
rect 4447 5179 4481 5195
rect 4447 4387 4481 4403
rect 4705 5179 4739 5195
rect 4705 4387 4739 4403
rect 4963 5179 4997 5195
rect 4963 4387 4997 4403
rect 5221 5179 5255 5195
rect 5221 4387 5255 4403
rect 5479 5179 5513 5195
rect 5479 4387 5513 4403
rect 5737 5179 5771 5195
rect 5737 4387 5771 4403
rect 5995 5179 6029 5195
rect 5995 4387 6029 4403
rect 6253 5179 6287 5195
rect 6253 4387 6287 4403
rect 6511 5179 6545 5195
rect 6511 4387 6545 4403
rect 81 4210 100 4358
rect 154 4210 173 4358
rect 365 4319 381 4353
rect 549 4319 565 4353
rect 623 4319 639 4353
rect 807 4319 823 4353
rect 881 4319 897 4353
rect 1065 4319 1081 4353
rect 1139 4319 1155 4353
rect 1323 4319 1339 4353
rect 1397 4319 1413 4353
rect 1581 4319 1597 4353
rect 1655 4319 1671 4353
rect 1839 4319 1855 4353
rect 1913 4319 1929 4353
rect 2097 4319 2113 4353
rect 2171 4319 2187 4353
rect 2355 4319 2371 4353
rect 2429 4319 2445 4353
rect 2613 4319 2629 4353
rect 2687 4319 2703 4353
rect 2871 4319 2887 4353
rect 2945 4319 2961 4353
rect 3129 4319 3145 4353
rect 3203 4319 3219 4353
rect 3387 4319 3403 4353
rect 3461 4319 3477 4353
rect 3645 4319 3661 4353
rect 3719 4319 3735 4353
rect 3903 4319 3919 4353
rect 3977 4319 3993 4353
rect 4161 4319 4177 4353
rect 4235 4319 4251 4353
rect 4419 4319 4435 4353
rect 4493 4319 4509 4353
rect 4677 4319 4693 4353
rect 4751 4319 4767 4353
rect 4935 4319 4951 4353
rect 5009 4319 5025 4353
rect 5193 4319 5209 4353
rect 5267 4319 5283 4353
rect 5451 4319 5467 4353
rect 5525 4319 5541 4353
rect 5709 4319 5725 4353
rect 5783 4319 5799 4353
rect 5967 4319 5983 4353
rect 6041 4319 6057 4353
rect 6225 4319 6241 4353
rect 6299 4319 6315 4353
rect 6483 4319 6499 4353
rect 81 2698 113 4210
rect 147 2708 173 4210
rect 365 3748 381 3782
rect 549 3748 565 3782
rect 623 3748 639 3782
rect 807 3748 823 3782
rect 881 3748 897 3782
rect 1065 3748 1081 3782
rect 1139 3748 1155 3782
rect 1323 3748 1339 3782
rect 1397 3748 1413 3782
rect 1581 3748 1597 3782
rect 1655 3748 1671 3782
rect 1839 3748 1855 3782
rect 1913 3748 1929 3782
rect 2097 3748 2113 3782
rect 2171 3748 2187 3782
rect 2355 3748 2371 3782
rect 2429 3748 2445 3782
rect 2613 3748 2629 3782
rect 2687 3748 2703 3782
rect 2871 3748 2887 3782
rect 2945 3748 2961 3782
rect 3129 3748 3145 3782
rect 3203 3748 3219 3782
rect 3387 3748 3403 3782
rect 3461 3748 3477 3782
rect 3645 3748 3661 3782
rect 3719 3748 3735 3782
rect 3903 3748 3919 3782
rect 3977 3748 3993 3782
rect 4161 3748 4177 3782
rect 4235 3748 4251 3782
rect 4419 3748 4435 3782
rect 4493 3748 4509 3782
rect 4677 3748 4693 3782
rect 4751 3748 4767 3782
rect 4935 3748 4951 3782
rect 5009 3748 5025 3782
rect 5193 3748 5209 3782
rect 5267 3748 5283 3782
rect 5451 3748 5467 3782
rect 5525 3748 5541 3782
rect 5709 3748 5725 3782
rect 5783 3748 5799 3782
rect 5967 3748 5983 3782
rect 6041 3748 6057 3782
rect 6225 3748 6241 3782
rect 6299 3748 6315 3782
rect 6483 3748 6499 3782
rect 319 3698 353 3714
rect 319 2906 353 2922
rect 577 3698 611 3714
rect 577 2906 611 2922
rect 835 3698 869 3714
rect 835 2906 869 2922
rect 1093 3698 1127 3714
rect 1093 2906 1127 2922
rect 1351 3698 1385 3714
rect 1351 2906 1385 2922
rect 1609 3698 1643 3714
rect 1609 2906 1643 2922
rect 1867 3698 1901 3714
rect 1867 2906 1901 2922
rect 2125 3698 2159 3714
rect 2125 2906 2159 2922
rect 2383 3698 2417 3714
rect 2383 2906 2417 2922
rect 2641 3698 2675 3714
rect 2641 2906 2675 2922
rect 2899 3698 2933 3714
rect 2899 2906 2933 2922
rect 3157 3698 3191 3714
rect 3157 2906 3191 2922
rect 3415 3698 3449 3714
rect 3415 2906 3449 2922
rect 3673 3698 3707 3714
rect 3673 2906 3707 2922
rect 3931 3698 3965 3714
rect 3931 2906 3965 2922
rect 4189 3698 4223 3714
rect 4189 2906 4223 2922
rect 4447 3698 4481 3714
rect 4447 2906 4481 2922
rect 4705 3698 4739 3714
rect 4705 2906 4739 2922
rect 4963 3698 4997 3714
rect 4963 2906 4997 2922
rect 5221 3698 5255 3714
rect 5221 2906 5255 2922
rect 5479 3698 5513 3714
rect 5479 2906 5513 2922
rect 5737 3698 5771 3714
rect 5737 2906 5771 2922
rect 5995 3698 6029 3714
rect 5995 2906 6029 2922
rect 6253 3698 6287 3714
rect 6253 2906 6287 2922
rect 6511 3698 6545 3714
rect 6511 2906 6545 2922
rect 365 2838 381 2872
rect 549 2838 565 2872
rect 623 2838 639 2872
rect 807 2838 823 2872
rect 881 2838 897 2872
rect 1065 2838 1081 2872
rect 1139 2838 1155 2872
rect 1323 2838 1339 2872
rect 1397 2838 1413 2872
rect 1581 2838 1597 2872
rect 1655 2838 1671 2872
rect 1839 2838 1855 2872
rect 1913 2838 1929 2872
rect 2097 2838 2113 2872
rect 2171 2838 2187 2872
rect 2355 2838 2371 2872
rect 2429 2838 2445 2872
rect 2613 2838 2629 2872
rect 2687 2838 2703 2872
rect 2871 2838 2887 2872
rect 2945 2838 2961 2872
rect 3129 2838 3145 2872
rect 3203 2838 3219 2872
rect 3387 2838 3403 2872
rect 3461 2838 3477 2872
rect 3645 2838 3661 2872
rect 3719 2838 3735 2872
rect 3903 2838 3919 2872
rect 3977 2838 3993 2872
rect 4161 2838 4177 2872
rect 4235 2838 4251 2872
rect 4419 2838 4435 2872
rect 4493 2838 4509 2872
rect 4677 2838 4693 2872
rect 4751 2838 4767 2872
rect 4935 2838 4951 2872
rect 5009 2838 5025 2872
rect 5193 2838 5209 2872
rect 5267 2838 5283 2872
rect 5451 2838 5467 2872
rect 5525 2838 5541 2872
rect 5709 2838 5725 2872
rect 5783 2838 5799 2872
rect 5967 2838 5983 2872
rect 6041 2838 6057 2872
rect 6225 2838 6241 2872
rect 6299 2838 6315 2872
rect 6483 2838 6499 2872
rect 6596 2715 6655 5321
rect 333 2708 6655 2715
rect 147 2698 6655 2708
rect 6689 2698 6712 5407
rect 81 2672 6712 2698
rect 81 2638 173 2672
rect 6629 2663 6712 2672
rect 81 2551 290 2638
rect 6631 2551 6712 2663
rect 81 2507 6712 2551
rect 80 2502 6712 2507
rect 80 2421 282 2502
rect 79 2406 282 2421
rect 809 2415 6712 2502
rect 809 2406 1367 2415
rect 79 2386 1367 2406
rect 79 2363 209 2386
rect 79 2329 113 2363
rect 147 2352 209 2363
rect 243 2352 299 2386
rect 333 2352 389 2386
rect 423 2352 479 2386
rect 513 2352 569 2386
rect 603 2352 659 2386
rect 693 2352 749 2386
rect 783 2352 839 2386
rect 873 2352 929 2386
rect 963 2352 1019 2386
rect 1053 2352 1109 2386
rect 1143 2352 1199 2386
rect 1233 2363 1367 2386
rect 1233 2352 1300 2363
rect 147 2329 1300 2352
rect 1334 2329 1367 2363
rect 79 2323 1367 2329
rect 79 2273 1183 2323
rect 79 2239 113 2273
rect 147 2239 1183 2273
rect 79 2205 373 2239
rect 407 2205 463 2239
rect 497 2205 553 2239
rect 587 2205 643 2239
rect 677 2205 733 2239
rect 767 2205 823 2239
rect 857 2205 913 2239
rect 947 2205 1003 2239
rect 1037 2205 1093 2239
rect 1127 2205 1183 2239
rect 79 2186 1183 2205
rect 79 2183 314 2186
rect 79 2149 113 2183
rect 147 2182 314 2183
rect 147 2149 261 2182
rect 79 2148 261 2149
rect 295 2148 314 2182
rect 79 2093 314 2148
rect 1132 2163 1183 2186
rect 1291 2273 1367 2323
rect 1291 2239 1300 2273
rect 1334 2239 1367 2273
rect 1291 2183 1367 2239
rect 1132 2129 1151 2163
rect 1291 2149 1300 2183
rect 1334 2149 1367 2183
rect 79 2059 113 2093
rect 147 2092 314 2093
rect 147 2059 261 2092
rect 79 2058 261 2059
rect 295 2058 314 2092
rect 79 2003 314 2058
rect 79 1969 113 2003
rect 147 2002 314 2003
rect 147 1969 261 2002
rect 79 1968 261 1969
rect 295 1968 314 2002
rect 79 1913 314 1968
rect 79 1879 113 1913
rect 147 1912 314 1913
rect 147 1890 261 1912
rect 79 1823 136 1879
rect 256 1878 261 1890
rect 295 1878 314 1912
rect 79 1789 113 1823
rect 256 1822 314 1878
rect 79 1733 136 1789
rect 256 1788 261 1822
rect 295 1788 314 1822
rect 79 1699 113 1733
rect 256 1732 314 1788
rect 79 1643 136 1699
rect 256 1698 261 1732
rect 295 1698 314 1732
rect 79 1609 113 1643
rect 256 1642 314 1698
rect 79 1553 136 1609
rect 256 1608 261 1642
rect 295 1608 314 1642
rect 79 1519 113 1553
rect 256 1552 314 1608
rect 79 1463 136 1519
rect 256 1518 261 1552
rect 295 1518 314 1552
rect 79 1429 113 1463
rect 256 1462 314 1518
rect 79 1411 136 1429
rect 256 1428 261 1462
rect 295 1428 314 1462
rect 376 2065 1070 2124
rect 376 2031 437 2065
rect 471 2037 527 2065
rect 561 2037 617 2065
rect 651 2037 707 2065
rect 483 2031 527 2037
rect 583 2031 617 2037
rect 683 2031 707 2037
rect 741 2037 797 2065
rect 741 2031 749 2037
rect 376 2003 449 2031
rect 483 2003 549 2031
rect 583 2003 649 2031
rect 683 2003 749 2031
rect 783 2031 797 2037
rect 831 2037 887 2065
rect 831 2031 849 2037
rect 783 2003 849 2031
rect 883 2031 887 2037
rect 921 2037 977 2065
rect 921 2031 949 2037
rect 1011 2031 1070 2065
rect 883 2003 949 2031
rect 983 2003 1070 2031
rect 376 1975 1070 2003
rect 376 1941 437 1975
rect 471 1941 527 1975
rect 561 1941 617 1975
rect 651 1941 707 1975
rect 741 1941 797 1975
rect 831 1941 887 1975
rect 921 1941 977 1975
rect 1011 1941 1070 1975
rect 376 1937 1070 1941
rect 376 1903 449 1937
rect 483 1903 549 1937
rect 583 1903 649 1937
rect 683 1903 749 1937
rect 783 1903 849 1937
rect 883 1903 949 1937
rect 983 1903 1070 1937
rect 376 1885 1070 1903
rect 376 1851 437 1885
rect 471 1851 527 1885
rect 561 1851 617 1885
rect 651 1851 707 1885
rect 741 1851 797 1885
rect 831 1851 887 1885
rect 921 1851 977 1885
rect 1011 1851 1070 1885
rect 376 1837 1070 1851
rect 376 1803 449 1837
rect 483 1803 549 1837
rect 583 1803 649 1837
rect 683 1803 749 1837
rect 783 1803 849 1837
rect 883 1803 949 1837
rect 983 1803 1070 1837
rect 376 1795 1070 1803
rect 376 1761 437 1795
rect 471 1761 527 1795
rect 561 1761 617 1795
rect 651 1761 707 1795
rect 741 1761 797 1795
rect 831 1761 887 1795
rect 921 1761 977 1795
rect 1011 1761 1070 1795
rect 376 1737 1070 1761
rect 376 1705 449 1737
rect 483 1705 549 1737
rect 583 1705 649 1737
rect 683 1705 749 1737
rect 376 1671 437 1705
rect 483 1703 527 1705
rect 583 1703 617 1705
rect 683 1703 707 1705
rect 471 1671 527 1703
rect 561 1671 617 1703
rect 651 1671 707 1703
rect 741 1703 749 1705
rect 783 1705 849 1737
rect 783 1703 797 1705
rect 741 1671 797 1703
rect 831 1703 849 1705
rect 883 1705 949 1737
rect 983 1705 1070 1737
rect 883 1703 887 1705
rect 831 1671 887 1703
rect 921 1703 949 1705
rect 921 1671 977 1703
rect 1011 1671 1070 1705
rect 376 1637 1070 1671
rect 376 1615 449 1637
rect 483 1615 549 1637
rect 583 1615 649 1637
rect 683 1615 749 1637
rect 376 1581 437 1615
rect 483 1603 527 1615
rect 583 1603 617 1615
rect 683 1603 707 1615
rect 471 1581 527 1603
rect 561 1581 617 1603
rect 651 1581 707 1603
rect 741 1603 749 1615
rect 783 1615 849 1637
rect 783 1603 797 1615
rect 741 1581 797 1603
rect 831 1603 849 1615
rect 883 1615 949 1637
rect 983 1615 1070 1637
rect 883 1603 887 1615
rect 831 1581 887 1603
rect 921 1603 949 1615
rect 921 1581 977 1603
rect 1011 1581 1070 1615
rect 376 1537 1070 1581
rect 376 1525 449 1537
rect 483 1525 549 1537
rect 583 1525 649 1537
rect 683 1525 749 1537
rect 376 1491 437 1525
rect 483 1503 527 1525
rect 583 1503 617 1525
rect 683 1503 707 1525
rect 471 1491 527 1503
rect 561 1491 617 1503
rect 651 1491 707 1503
rect 741 1503 749 1525
rect 783 1525 849 1537
rect 783 1503 797 1525
rect 741 1491 797 1503
rect 831 1503 849 1525
rect 883 1525 949 1537
rect 983 1525 1070 1537
rect 883 1503 887 1525
rect 831 1491 887 1503
rect 921 1503 949 1525
rect 921 1491 977 1503
rect 1011 1491 1070 1525
rect 376 1430 1070 1491
rect 1132 2073 1183 2129
rect 1291 2093 1367 2149
rect 1132 2039 1151 2073
rect 1291 2059 1300 2093
rect 1334 2059 1367 2093
rect 1132 1983 1183 2039
rect 1291 2003 1367 2059
rect 1132 1949 1151 1983
rect 1291 1969 1300 2003
rect 1334 1969 1367 2003
rect 1132 1893 1183 1949
rect 1291 1913 1367 1969
rect 1990 1950 6712 2415
rect 1990 1941 7613 1950
rect 1132 1859 1151 1893
rect 1291 1879 1300 1913
rect 1334 1879 1367 1913
rect 1132 1803 1183 1859
rect 1291 1823 1367 1879
rect 1132 1769 1151 1803
rect 1291 1789 1300 1823
rect 1334 1789 1367 1823
rect 1132 1713 1183 1769
rect 1291 1733 1367 1789
rect 1132 1679 1151 1713
rect 1291 1699 1300 1733
rect 1334 1699 1367 1733
rect 1132 1623 1183 1679
rect 1291 1643 1367 1699
rect 1132 1589 1151 1623
rect 1291 1609 1300 1643
rect 1334 1609 1367 1643
rect 1132 1533 1183 1589
rect 1291 1553 1367 1609
rect 1132 1499 1151 1533
rect 1291 1519 1300 1553
rect 1334 1519 1367 1553
rect 1132 1443 1183 1499
rect 1291 1463 1367 1519
rect 256 1411 314 1428
rect 79 1373 314 1411
rect 79 1339 113 1373
rect 147 1368 314 1373
rect 1132 1409 1151 1443
rect 1291 1429 1300 1463
rect 1334 1429 1367 1463
rect 1132 1368 1183 1409
rect 147 1349 1183 1368
rect 147 1339 339 1349
rect 79 1315 339 1339
rect 373 1315 429 1349
rect 463 1315 519 1349
rect 553 1315 609 1349
rect 643 1315 699 1349
rect 733 1315 789 1349
rect 823 1315 879 1349
rect 913 1315 969 1349
rect 1003 1315 1059 1349
rect 1093 1315 1183 1349
rect 79 1313 1183 1315
rect 79 1283 233 1313
rect 79 1249 113 1283
rect 147 1249 233 1283
rect 79 1199 233 1249
rect 1058 1280 1183 1313
rect 1291 1373 1367 1429
rect 1291 1339 1300 1373
rect 1334 1339 1367 1373
rect 1291 1283 1367 1339
rect 1291 1280 1300 1283
rect 1058 1249 1300 1280
rect 1334 1249 1367 1283
rect 1058 1199 1367 1249
rect 79 1165 209 1199
rect 1058 1165 1109 1199
rect 1143 1165 1199 1199
rect 1233 1165 1367 1199
rect 79 1133 1367 1165
rect 1991 1922 7613 1941
rect 1991 1760 2084 1922
rect 7491 1820 7613 1922
rect 7506 1786 7613 1820
rect 1991 1178 2038 1760
rect 2072 1731 2084 1760
rect 7491 1760 7613 1786
rect 7491 1731 7532 1760
rect 2072 1694 7532 1731
rect 2072 1199 2114 1694
rect 2251 1612 2267 1646
rect 2435 1612 2451 1646
rect 2509 1612 2525 1646
rect 2693 1612 2709 1646
rect 2767 1612 2783 1646
rect 2951 1612 2967 1646
rect 3025 1612 3041 1646
rect 3209 1612 3225 1646
rect 3283 1612 3299 1646
rect 3467 1612 3483 1646
rect 3541 1612 3557 1646
rect 3725 1612 3741 1646
rect 3799 1612 3815 1646
rect 3983 1612 3999 1646
rect 4057 1612 4073 1646
rect 4241 1612 4257 1646
rect 4315 1612 4331 1646
rect 4499 1612 4515 1646
rect 4573 1612 4589 1646
rect 4757 1612 4773 1646
rect 4831 1612 4847 1646
rect 5015 1612 5031 1646
rect 5089 1612 5105 1646
rect 5273 1612 5289 1646
rect 5347 1612 5363 1646
rect 5531 1612 5547 1646
rect 5605 1612 5621 1646
rect 5789 1612 5805 1646
rect 5863 1612 5879 1646
rect 6047 1612 6063 1646
rect 6121 1612 6137 1646
rect 6305 1612 6321 1646
rect 6379 1612 6395 1646
rect 6563 1612 6579 1646
rect 6637 1612 6653 1646
rect 6821 1612 6837 1646
rect 6895 1612 6911 1646
rect 7079 1612 7095 1646
rect 7153 1612 7169 1646
rect 7337 1612 7353 1646
rect 2205 1562 2239 1578
rect 2205 1370 2239 1386
rect 2463 1562 2497 1578
rect 2463 1370 2497 1386
rect 2721 1562 2755 1578
rect 2721 1370 2755 1386
rect 2979 1562 3013 1578
rect 2979 1370 3013 1386
rect 3237 1562 3271 1578
rect 3237 1370 3271 1386
rect 3495 1562 3529 1578
rect 3495 1370 3529 1386
rect 3753 1562 3787 1578
rect 3753 1370 3787 1386
rect 4011 1562 4045 1578
rect 4011 1370 4045 1386
rect 4269 1562 4303 1578
rect 4269 1370 4303 1386
rect 4527 1562 4561 1578
rect 4527 1370 4561 1386
rect 4785 1562 4819 1578
rect 4785 1370 4819 1386
rect 5043 1562 5077 1578
rect 5043 1370 5077 1386
rect 5301 1562 5335 1578
rect 5301 1370 5335 1386
rect 5559 1562 5593 1578
rect 5559 1370 5593 1386
rect 5817 1562 5851 1578
rect 5817 1370 5851 1386
rect 6075 1562 6109 1578
rect 6075 1370 6109 1386
rect 6333 1562 6367 1578
rect 6333 1370 6367 1386
rect 6591 1562 6625 1578
rect 6591 1370 6625 1386
rect 6849 1562 6883 1578
rect 6849 1370 6883 1386
rect 7107 1562 7141 1578
rect 7107 1370 7141 1386
rect 7365 1562 7399 1578
rect 7365 1370 7399 1386
rect 2251 1302 2267 1336
rect 2435 1302 2451 1336
rect 2509 1302 2525 1336
rect 2693 1302 2709 1336
rect 2767 1302 2783 1336
rect 2951 1302 2967 1336
rect 3025 1302 3041 1336
rect 3209 1302 3225 1336
rect 3283 1302 3299 1336
rect 3467 1302 3483 1336
rect 3541 1302 3557 1336
rect 3725 1302 3741 1336
rect 3799 1302 3815 1336
rect 3983 1302 3999 1336
rect 4057 1302 4073 1336
rect 4241 1302 4257 1336
rect 4315 1302 4331 1336
rect 4499 1302 4515 1336
rect 4573 1302 4589 1336
rect 4757 1302 4773 1336
rect 4831 1302 4847 1336
rect 5015 1302 5031 1336
rect 5089 1302 5105 1336
rect 5273 1302 5289 1336
rect 5347 1302 5363 1336
rect 5531 1302 5547 1336
rect 5605 1302 5621 1336
rect 5789 1302 5805 1336
rect 5863 1302 5879 1336
rect 6047 1302 6063 1336
rect 6121 1302 6137 1336
rect 6305 1302 6321 1336
rect 6379 1302 6395 1336
rect 6563 1302 6579 1336
rect 6637 1302 6653 1336
rect 6821 1302 6837 1336
rect 6895 1302 6911 1336
rect 7079 1302 7095 1336
rect 7153 1302 7169 1336
rect 7337 1302 7353 1336
rect 7490 1199 7532 1694
rect 2072 1178 7532 1199
rect 7566 1178 7613 1760
rect 1991 1152 7613 1178
rect 1991 1118 2098 1152
rect 7506 1118 7613 1152
rect 1991 1060 7613 1118
rect 2386 990 3153 992
rect 2384 970 3153 990
rect 51 912 239 960
rect 1347 912 1604 960
rect 1881 912 1992 960
rect 51 793 103 912
rect 1943 877 1992 912
rect 247 833 263 867
rect 631 833 647 867
rect 705 833 721 867
rect 1089 833 1105 867
rect 1372 833 1388 867
rect 1556 833 1572 867
rect 1630 833 1646 867
rect 1814 833 1830 867
rect 201 774 235 790
rect 201 682 235 698
rect 659 774 693 790
rect 659 682 693 698
rect 1117 774 1151 790
rect 1117 682 1151 698
rect 1326 774 1360 790
rect 247 605 263 639
rect 631 605 647 639
rect 705 605 721 639
rect 1089 605 1105 639
rect 1326 582 1360 598
rect 1584 774 1618 790
rect 1584 582 1618 598
rect 1842 774 1876 790
rect 1842 582 1876 598
rect 51 468 103 557
rect 1372 505 1388 539
rect 1556 505 1572 539
rect 1630 505 1646 539
rect 1814 505 1830 539
rect 1911 498 1943 531
rect 2384 936 2503 970
rect 3031 936 3153 970
rect 2384 924 3153 936
rect 3663 970 4453 986
rect 3663 936 3793 970
rect 4321 936 4453 970
rect 2384 874 2462 924
rect 2384 531 2407 874
rect 1992 500 2407 531
rect 2441 531 2462 874
rect 3074 874 3152 924
rect 3663 910 4453 936
rect 2567 834 2583 868
rect 2951 834 2967 868
rect 2521 775 2555 791
rect 2521 583 2555 599
rect 2979 775 3013 791
rect 2979 583 3013 599
rect 2441 500 2465 531
rect 2567 506 2583 540
rect 2951 506 2967 540
rect 1992 498 2465 500
rect -26 467 214 468
rect 260 467 1248 468
rect -26 465 1248 467
rect 1911 465 2465 498
rect -26 462 2465 465
rect -26 439 199 462
rect 1874 458 2465 462
rect 3074 500 3093 874
rect 3127 808 3152 874
rect 3667 874 3752 910
rect 3667 808 3697 874
rect 3127 500 3697 808
rect 3731 500 3752 874
rect 4373 874 4453 910
rect 3857 834 3873 868
rect 4241 834 4257 868
rect 3811 775 3845 791
rect 3811 583 3845 599
rect 4269 775 4303 791
rect 4269 583 4303 599
rect 3857 506 3873 540
rect 4241 506 4257 540
rect 3074 458 3752 500
rect 4373 500 4383 874
rect 4417 820 4453 874
rect 4959 970 5743 995
rect 6253 984 7623 986
rect 4959 936 5083 970
rect 5611 936 5743 970
rect 4959 912 5743 936
rect 4959 874 5050 912
rect 4959 820 4987 874
rect 4417 500 4987 820
rect 5021 500 5050 874
rect 5647 874 5743 912
rect 5147 834 5163 868
rect 5531 834 5547 868
rect 5101 775 5135 791
rect 5101 583 5135 599
rect 5559 775 5593 791
rect 5559 583 5593 599
rect 5147 506 5163 540
rect 5531 506 5547 540
rect 4373 459 5050 500
rect 5647 500 5673 874
rect 5707 820 5743 874
rect 6251 946 7623 984
rect 6251 912 6350 946
rect 7514 912 7623 946
rect 6251 907 7623 912
rect 6251 886 6336 907
rect 6251 820 6290 886
rect 5707 500 6290 820
rect 5647 462 6290 500
rect 6324 462 6336 886
rect 7519 886 7623 907
rect 6437 834 6453 868
rect 6821 834 6837 868
rect 7018 834 7034 868
rect 7402 834 7418 868
rect 6391 775 6425 791
rect 6391 583 6425 599
rect 6849 775 6883 791
rect 6849 583 6883 599
rect 6972 775 7006 791
rect 6972 583 7006 599
rect 7430 775 7464 791
rect 7430 583 7464 599
rect 6437 506 6453 540
rect 6821 506 6837 540
rect 7018 506 7034 540
rect 7402 506 7418 540
rect 5647 459 6336 462
rect 4373 458 5146 459
rect 5646 458 6336 459
rect 7519 462 7540 886
rect 7574 462 7623 886
rect 7519 458 7623 462
rect 1874 442 7623 458
rect 1874 441 7622 442
rect -26 307 24 439
rect 1916 438 7622 441
rect 1916 406 2503 438
rect 2003 404 2503 406
rect 3031 404 3793 438
rect 4321 404 5083 438
rect 5611 436 7622 438
rect 5611 404 6350 436
rect 2003 402 6350 404
rect 7514 402 7622 436
rect 2003 328 7622 402
rect -26 306 1017 307
rect 2003 306 2514 328
rect -26 228 2514 306
rect -26 80 25 228
rect 2004 189 2514 228
rect 7509 189 7622 328
rect 2004 158 7622 189
rect 2004 80 7629 158
rect -26 34 7629 80
rect -25 0 7629 34
rect -25 -2 2035 0
<< viali >>
rect 97 5467 6675 5604
rect 97 5433 173 5467
rect 173 5433 6629 5467
rect 6629 5433 6675 5467
rect 97 5430 6675 5433
rect 100 5196 113 5348
rect 113 5196 147 5348
rect 147 5196 154 5348
rect 381 5229 549 5263
rect 639 5229 807 5263
rect 897 5229 1065 5263
rect 1155 5229 1323 5263
rect 1413 5229 1581 5263
rect 1671 5229 1839 5263
rect 1929 5229 2097 5263
rect 2187 5229 2355 5263
rect 2445 5229 2613 5263
rect 2703 5229 2871 5263
rect 2961 5229 3129 5263
rect 3219 5229 3387 5263
rect 3477 5229 3645 5263
rect 3735 5229 3903 5263
rect 3993 5229 4161 5263
rect 4251 5229 4419 5263
rect 4509 5229 4677 5263
rect 4767 5229 4935 5263
rect 5025 5229 5193 5263
rect 5283 5229 5451 5263
rect 5541 5229 5709 5263
rect 5799 5229 5967 5263
rect 6057 5229 6225 5263
rect 6315 5229 6483 5263
rect 319 4403 353 5179
rect 577 4403 611 5179
rect 835 4403 869 5179
rect 1093 4403 1127 5179
rect 1351 4403 1385 5179
rect 1609 4403 1643 5179
rect 1867 4403 1901 5179
rect 2125 4403 2159 5179
rect 2383 4403 2417 5179
rect 2641 4403 2675 5179
rect 2899 4403 2933 5179
rect 3157 4403 3191 5179
rect 3415 4403 3449 5179
rect 3673 4403 3707 5179
rect 3931 4403 3965 5179
rect 4189 4403 4223 5179
rect 4447 4403 4481 5179
rect 4705 4403 4739 5179
rect 4963 4403 4997 5179
rect 5221 4403 5255 5179
rect 5479 4403 5513 5179
rect 5737 4403 5771 5179
rect 5995 4403 6029 5179
rect 6253 4403 6287 5179
rect 6511 4403 6545 5179
rect 100 4210 113 4358
rect 113 4210 147 4358
rect 147 4210 154 4358
rect 381 4319 549 4353
rect 639 4319 807 4353
rect 897 4319 1065 4353
rect 1155 4319 1323 4353
rect 1413 4319 1581 4353
rect 1671 4319 1839 4353
rect 1929 4319 2097 4353
rect 2187 4319 2355 4353
rect 2445 4319 2613 4353
rect 2703 4319 2871 4353
rect 2961 4319 3129 4353
rect 3219 4319 3387 4353
rect 3477 4319 3645 4353
rect 3735 4319 3903 4353
rect 3993 4319 4161 4353
rect 4251 4319 4419 4353
rect 4509 4319 4677 4353
rect 4767 4319 4935 4353
rect 5025 4319 5193 4353
rect 5283 4319 5451 4353
rect 5541 4319 5709 4353
rect 5799 4319 5967 4353
rect 6057 4319 6225 4353
rect 6315 4319 6483 4353
rect 381 3748 549 3782
rect 639 3748 807 3782
rect 897 3748 1065 3782
rect 1155 3748 1323 3782
rect 1413 3748 1581 3782
rect 1671 3748 1839 3782
rect 1929 3748 2097 3782
rect 2187 3748 2355 3782
rect 2445 3748 2613 3782
rect 2703 3748 2871 3782
rect 2961 3748 3129 3782
rect 3219 3748 3387 3782
rect 3477 3748 3645 3782
rect 3735 3748 3903 3782
rect 3993 3748 4161 3782
rect 4251 3748 4419 3782
rect 4509 3748 4677 3782
rect 4767 3748 4935 3782
rect 5025 3748 5193 3782
rect 5283 3748 5451 3782
rect 5541 3748 5709 3782
rect 5799 3748 5967 3782
rect 6057 3748 6225 3782
rect 6315 3748 6483 3782
rect 319 2922 353 3698
rect 577 2922 611 3698
rect 835 2922 869 3698
rect 1093 2922 1127 3698
rect 1351 2922 1385 3698
rect 1609 2922 1643 3698
rect 1867 2922 1901 3698
rect 2125 2922 2159 3698
rect 2383 2922 2417 3698
rect 2641 2922 2675 3698
rect 2899 2922 2933 3698
rect 3157 2922 3191 3698
rect 3415 2922 3449 3698
rect 3673 2922 3707 3698
rect 3931 2922 3965 3698
rect 4189 2922 4223 3698
rect 4447 2922 4481 3698
rect 4705 2922 4739 3698
rect 4963 2922 4997 3698
rect 5221 2922 5255 3698
rect 5479 2922 5513 3698
rect 5737 2922 5771 3698
rect 5995 2922 6029 3698
rect 6253 2922 6287 3698
rect 6511 2922 6545 3698
rect 381 2838 549 2872
rect 639 2838 807 2872
rect 897 2838 1065 2872
rect 1155 2838 1323 2872
rect 1413 2838 1581 2872
rect 1671 2838 1839 2872
rect 1929 2838 2097 2872
rect 2187 2838 2355 2872
rect 2445 2838 2613 2872
rect 2703 2838 2871 2872
rect 2961 2838 3129 2872
rect 3219 2838 3387 2872
rect 3477 2838 3645 2872
rect 3735 2838 3903 2872
rect 3993 2838 4161 2872
rect 4251 2838 4419 2872
rect 4509 2838 4677 2872
rect 4767 2838 4935 2872
rect 5025 2838 5193 2872
rect 5283 2838 5451 2872
rect 5541 2838 5709 2872
rect 5799 2838 5967 2872
rect 6057 2838 6225 2872
rect 6315 2838 6483 2872
rect 290 2638 6629 2663
rect 6629 2638 6631 2663
rect 290 2551 6631 2638
rect 282 2406 809 2502
rect 1183 2163 1291 2323
rect 1183 2129 1185 2163
rect 1185 2129 1291 2163
rect 136 1879 147 1890
rect 147 1879 256 1890
rect 136 1823 256 1879
rect 136 1789 147 1823
rect 147 1789 256 1823
rect 136 1733 256 1789
rect 136 1699 147 1733
rect 147 1699 256 1733
rect 136 1643 256 1699
rect 136 1609 147 1643
rect 147 1609 256 1643
rect 136 1553 256 1609
rect 136 1519 147 1553
rect 147 1519 256 1553
rect 136 1463 256 1519
rect 136 1429 147 1463
rect 147 1429 256 1463
rect 136 1411 256 1429
rect 449 2031 471 2037
rect 471 2031 483 2037
rect 549 2031 561 2037
rect 561 2031 583 2037
rect 649 2031 651 2037
rect 651 2031 683 2037
rect 449 2003 483 2031
rect 549 2003 583 2031
rect 649 2003 683 2031
rect 749 2003 783 2037
rect 849 2003 883 2037
rect 949 2031 977 2037
rect 977 2031 983 2037
rect 949 2003 983 2031
rect 449 1903 483 1937
rect 549 1903 583 1937
rect 649 1903 683 1937
rect 749 1903 783 1937
rect 849 1903 883 1937
rect 949 1903 983 1937
rect 449 1803 483 1837
rect 549 1803 583 1837
rect 649 1803 683 1837
rect 749 1803 783 1837
rect 849 1803 883 1837
rect 949 1803 983 1837
rect 449 1705 483 1737
rect 549 1705 583 1737
rect 649 1705 683 1737
rect 449 1703 471 1705
rect 471 1703 483 1705
rect 549 1703 561 1705
rect 561 1703 583 1705
rect 649 1703 651 1705
rect 651 1703 683 1705
rect 749 1703 783 1737
rect 849 1703 883 1737
rect 949 1705 983 1737
rect 949 1703 977 1705
rect 977 1703 983 1705
rect 449 1615 483 1637
rect 549 1615 583 1637
rect 649 1615 683 1637
rect 449 1603 471 1615
rect 471 1603 483 1615
rect 549 1603 561 1615
rect 561 1603 583 1615
rect 649 1603 651 1615
rect 651 1603 683 1615
rect 749 1603 783 1637
rect 849 1603 883 1637
rect 949 1615 983 1637
rect 949 1603 977 1615
rect 977 1603 983 1615
rect 449 1525 483 1537
rect 549 1525 583 1537
rect 649 1525 683 1537
rect 449 1503 471 1525
rect 471 1503 483 1525
rect 549 1503 561 1525
rect 561 1503 583 1525
rect 649 1503 651 1525
rect 651 1503 683 1525
rect 749 1503 783 1537
rect 849 1503 883 1537
rect 949 1525 983 1537
rect 949 1503 977 1525
rect 977 1503 983 1525
rect 1183 2073 1291 2129
rect 1183 2039 1185 2073
rect 1185 2039 1291 2073
rect 1183 1983 1291 2039
rect 1183 1949 1185 1983
rect 1185 1949 1291 1983
rect 1183 1893 1291 1949
rect 1183 1859 1185 1893
rect 1185 1859 1291 1893
rect 1183 1803 1291 1859
rect 1183 1769 1185 1803
rect 1185 1769 1291 1803
rect 1183 1713 1291 1769
rect 1183 1679 1185 1713
rect 1185 1679 1291 1713
rect 1183 1623 1291 1679
rect 1183 1589 1185 1623
rect 1185 1589 1291 1623
rect 1183 1533 1291 1589
rect 1183 1499 1185 1533
rect 1185 1499 1291 1533
rect 1183 1443 1291 1499
rect 1183 1409 1185 1443
rect 1185 1409 1291 1443
rect 233 1199 1058 1313
rect 1183 1280 1291 1409
rect 233 1165 243 1199
rect 243 1165 299 1199
rect 299 1165 333 1199
rect 333 1165 389 1199
rect 389 1165 423 1199
rect 423 1165 479 1199
rect 479 1165 513 1199
rect 513 1165 569 1199
rect 569 1165 603 1199
rect 603 1165 659 1199
rect 659 1165 693 1199
rect 693 1165 749 1199
rect 749 1165 783 1199
rect 783 1165 839 1199
rect 839 1165 873 1199
rect 873 1165 929 1199
rect 929 1165 963 1199
rect 963 1165 1019 1199
rect 1019 1165 1053 1199
rect 1053 1165 1058 1199
rect 2084 1820 7491 1922
rect 2084 1786 2098 1820
rect 2098 1786 7491 1820
rect 2084 1731 7491 1786
rect 2267 1612 2435 1646
rect 2525 1612 2693 1646
rect 2783 1612 2951 1646
rect 3041 1612 3209 1646
rect 3299 1612 3467 1646
rect 3557 1612 3725 1646
rect 3815 1612 3983 1646
rect 4073 1612 4241 1646
rect 4331 1612 4499 1646
rect 4589 1612 4757 1646
rect 4847 1612 5015 1646
rect 5105 1612 5273 1646
rect 5363 1612 5531 1646
rect 5621 1612 5789 1646
rect 5879 1612 6047 1646
rect 6137 1612 6305 1646
rect 6395 1612 6563 1646
rect 6653 1612 6821 1646
rect 6911 1612 7079 1646
rect 7169 1612 7337 1646
rect 2205 1386 2239 1562
rect 2463 1386 2497 1562
rect 2721 1386 2755 1562
rect 2979 1386 3013 1562
rect 3237 1386 3271 1562
rect 3495 1386 3529 1562
rect 3753 1386 3787 1562
rect 4011 1386 4045 1562
rect 4269 1386 4303 1562
rect 4527 1386 4561 1562
rect 4785 1386 4819 1562
rect 5043 1386 5077 1562
rect 5301 1386 5335 1562
rect 5559 1386 5593 1562
rect 5817 1386 5851 1562
rect 6075 1386 6109 1562
rect 6333 1386 6367 1562
rect 6591 1386 6625 1562
rect 6849 1386 6883 1562
rect 7107 1386 7141 1562
rect 7365 1386 7399 1562
rect 2267 1302 2435 1336
rect 2525 1302 2693 1336
rect 2783 1302 2951 1336
rect 3041 1302 3209 1336
rect 3299 1302 3467 1336
rect 3557 1302 3725 1336
rect 3815 1302 3983 1336
rect 4073 1302 4241 1336
rect 4331 1302 4499 1336
rect 4589 1302 4757 1336
rect 4847 1302 5015 1336
rect 5105 1302 5273 1336
rect 5363 1302 5531 1336
rect 5621 1302 5789 1336
rect 5879 1302 6047 1336
rect 6137 1302 6305 1336
rect 6395 1302 6563 1336
rect 6653 1302 6821 1336
rect 6911 1302 7079 1336
rect 7169 1302 7337 1336
rect 263 833 631 867
rect 721 833 1089 867
rect 1388 833 1556 867
rect 1646 833 1814 867
rect 201 698 235 774
rect 659 698 693 774
rect 1117 698 1151 774
rect 263 605 631 639
rect 721 605 1089 639
rect 1326 598 1360 774
rect 1584 598 1618 774
rect 1842 598 1876 774
rect 1388 505 1556 539
rect 1646 505 1814 539
rect 2583 834 2951 868
rect 2521 599 2555 775
rect 2979 599 3013 775
rect 2583 506 2951 540
rect 3873 834 4241 868
rect 3811 599 3845 775
rect 4269 599 4303 775
rect 3873 506 4241 540
rect 5163 834 5531 868
rect 5101 599 5135 775
rect 5559 599 5593 775
rect 5163 506 5531 540
rect 6453 834 6821 868
rect 7034 834 7402 868
rect 6391 599 6425 775
rect 6849 599 6883 775
rect 6972 599 7006 775
rect 7430 599 7464 775
rect 6453 506 6821 540
rect 7034 506 7402 540
rect 1017 439 1874 441
rect 24 410 199 439
rect 199 410 1874 439
rect 1874 410 1916 441
rect 24 406 1916 410
rect 24 307 2003 406
rect 1017 306 2003 307
rect 25 80 2004 228
rect 2514 189 7509 328
<< metal1 >>
rect 85 5604 6687 5610
rect 85 5430 97 5604
rect 6675 5430 6687 5604
rect 85 5424 6687 5430
rect 94 5348 160 5360
rect 90 5196 100 5348
rect 154 5196 164 5348
rect 369 5263 819 5269
rect 369 5229 381 5263
rect 549 5229 639 5263
rect 807 5229 819 5263
rect 369 5223 819 5229
rect 885 5263 1335 5269
rect 885 5229 897 5263
rect 1065 5229 1155 5263
rect 1323 5229 1335 5263
rect 885 5223 1335 5229
rect 1401 5263 2367 5269
rect 1401 5229 1413 5263
rect 1581 5229 1671 5263
rect 1839 5229 1929 5263
rect 2097 5229 2187 5263
rect 2355 5229 2367 5263
rect 1401 5223 2367 5229
rect 2433 5263 2883 5269
rect 2433 5229 2445 5263
rect 2613 5229 2703 5263
rect 2871 5229 2883 5263
rect 2433 5223 2883 5229
rect 2949 5263 3915 5269
rect 2949 5229 2961 5263
rect 3129 5229 3219 5263
rect 3387 5229 3477 5263
rect 3645 5229 3735 5263
rect 3903 5229 3915 5263
rect 2949 5223 3915 5229
rect 3981 5263 4431 5269
rect 3981 5229 3993 5263
rect 4161 5229 4251 5263
rect 4419 5229 4431 5263
rect 3981 5223 4431 5229
rect 4497 5263 5463 5269
rect 4497 5229 4509 5263
rect 4677 5229 4767 5263
rect 4935 5229 5025 5263
rect 5193 5229 5283 5263
rect 5451 5229 5463 5263
rect 4497 5223 5463 5229
rect 5529 5263 5979 5269
rect 5529 5229 5541 5263
rect 5709 5229 5799 5263
rect 5967 5229 5979 5263
rect 5529 5223 5979 5229
rect 6045 5263 6495 5269
rect 6045 5229 6057 5263
rect 6225 5229 6315 5263
rect 6483 5229 6495 5263
rect 6045 5223 6495 5229
rect 94 5184 160 5196
rect 313 5179 359 5191
rect 294 4979 304 5179
rect 368 4979 378 5179
rect 313 4403 319 4979
rect 353 4403 359 4979
rect 313 4391 359 4403
rect 94 4358 160 4370
rect 418 4359 507 5223
rect 571 5179 617 5191
rect 571 4603 577 5179
rect 611 4603 617 5179
rect 556 4403 566 4603
rect 622 4403 632 4603
rect 571 4391 617 4403
rect 682 4362 771 5223
rect 829 5179 875 5191
rect 829 4827 835 5179
rect 869 4827 875 5179
rect 931 4827 1020 5223
rect 1087 5179 1133 5191
rect 1074 4979 1084 5179
rect 1136 4979 1146 5179
rect 816 4727 826 4827
rect 878 4727 888 4827
rect 931 4727 950 4827
rect 1002 4727 1020 4827
rect 829 4403 835 4727
rect 869 4403 875 4727
rect 829 4391 875 4403
rect 682 4359 707 4362
rect 90 4210 100 4358
rect 154 4210 164 4358
rect 369 4353 707 4359
rect 807 4359 817 4362
rect 931 4359 1020 4727
rect 1087 4403 1093 4979
rect 1127 4403 1133 4979
rect 1087 4391 1133 4403
rect 1195 4827 1283 5223
rect 1345 5179 1391 5191
rect 1345 4827 1351 5179
rect 1385 4827 1391 5179
rect 1195 4727 1215 4827
rect 1267 4727 1283 4827
rect 1332 4727 1342 4827
rect 1394 4727 1404 4827
rect 1195 4362 1283 4727
rect 1345 4403 1351 4727
rect 1385 4403 1391 4727
rect 1345 4391 1391 4403
rect 1195 4359 1223 4362
rect 369 4319 381 4353
rect 549 4319 639 4353
rect 369 4313 707 4319
rect 697 4310 707 4313
rect 807 4313 819 4359
rect 885 4353 1223 4359
rect 1323 4359 1333 4362
rect 1456 4359 1544 5223
rect 1603 5179 1649 5191
rect 1603 4603 1609 5179
rect 1643 4603 1649 5179
rect 1588 4403 1598 4603
rect 1654 4403 1664 4603
rect 1603 4391 1649 4403
rect 1719 4359 1807 5223
rect 1861 5179 1907 5191
rect 1842 4979 1852 5179
rect 1916 4979 1926 5179
rect 1861 4403 1867 4979
rect 1901 4403 1907 4979
rect 1861 4391 1907 4403
rect 1969 4359 2057 5223
rect 2119 5179 2165 5191
rect 2119 4603 2125 5179
rect 2159 4603 2165 5179
rect 2104 4403 2114 4603
rect 2170 4403 2180 4603
rect 2119 4391 2165 4403
rect 2228 4372 2316 5223
rect 2377 5179 2423 5191
rect 2377 4827 2383 5179
rect 2417 4827 2423 5179
rect 2481 4828 2574 5223
rect 2635 5179 2681 5191
rect 2622 4979 2632 5179
rect 2684 4979 2694 5179
rect 2364 4727 2374 4827
rect 2426 4727 2436 4827
rect 2481 4728 2497 4828
rect 2549 4728 2574 4828
rect 2377 4403 2383 4727
rect 2417 4403 2423 4727
rect 2377 4391 2423 4403
rect 2206 4362 2316 4372
rect 2206 4359 2229 4362
rect 885 4319 897 4353
rect 1065 4319 1155 4353
rect 885 4313 1223 4319
rect 807 4310 817 4313
rect 1213 4310 1223 4313
rect 1323 4313 1335 4359
rect 1401 4353 2229 4359
rect 2355 4359 2365 4362
rect 2481 4359 2574 4728
rect 2635 4403 2641 4979
rect 2675 4403 2681 4979
rect 2635 4391 2681 4403
rect 2743 4826 2831 5223
rect 2893 5179 2939 5191
rect 2893 4827 2899 5179
rect 2933 4827 2939 5179
rect 2743 4726 2759 4826
rect 2811 4726 2831 4826
rect 2880 4727 2890 4827
rect 2942 4727 2952 4827
rect 2743 4362 2831 4726
rect 2893 4403 2899 4727
rect 2933 4403 2939 4727
rect 2893 4391 2939 4403
rect 2743 4359 2771 4362
rect 1401 4319 1413 4353
rect 1581 4319 1671 4353
rect 1839 4319 1929 4353
rect 2097 4319 2187 4353
rect 1401 4313 2229 4319
rect 1323 4310 1333 4313
rect 2206 4310 2229 4313
rect 2355 4313 2367 4359
rect 2433 4353 2771 4359
rect 2871 4359 2881 4362
rect 3008 4359 3096 5223
rect 3151 5179 3197 5191
rect 3151 4603 3157 5179
rect 3191 4603 3197 5179
rect 3136 4403 3146 4603
rect 3202 4403 3212 4603
rect 3151 4391 3197 4403
rect 3264 4359 3352 5223
rect 3409 5179 3455 5191
rect 3390 4979 3400 5179
rect 3464 4979 3474 5179
rect 3409 4403 3415 4979
rect 3449 4403 3455 4979
rect 3409 4391 3455 4403
rect 3521 4359 3609 5223
rect 3667 5179 3713 5191
rect 3667 4603 3673 5179
rect 3707 4603 3713 5179
rect 3652 4403 3662 4603
rect 3718 4403 3728 4603
rect 3667 4391 3713 4403
rect 3780 4362 3868 5223
rect 3925 5179 3971 5191
rect 3925 4827 3931 5179
rect 3965 4827 3971 5179
rect 3912 4727 3922 4827
rect 3974 4727 3984 4827
rect 4032 4825 4120 5223
rect 4183 5179 4229 5191
rect 4169 4979 4179 5179
rect 4231 4979 4241 5179
rect 3925 4403 3931 4727
rect 3965 4403 3971 4727
rect 3925 4391 3971 4403
rect 4032 4725 4052 4825
rect 4104 4725 4120 4825
rect 3763 4359 3777 4362
rect 2433 4319 2445 4353
rect 2613 4319 2703 4353
rect 2433 4313 2771 4319
rect 2355 4310 2365 4313
rect 2761 4310 2771 4313
rect 2871 4313 2883 4359
rect 2949 4353 3777 4359
rect 3903 4359 3913 4362
rect 4032 4359 4120 4725
rect 4183 4403 4189 4979
rect 4223 4403 4229 4979
rect 4183 4391 4229 4403
rect 4289 4828 4377 5223
rect 4289 4728 4304 4828
rect 4356 4728 4377 4828
rect 4441 5179 4487 5191
rect 4441 4827 4447 5179
rect 4481 4827 4487 5179
rect 4289 4362 4377 4728
rect 4428 4727 4438 4827
rect 4490 4727 4500 4827
rect 4441 4403 4447 4727
rect 4481 4403 4487 4727
rect 4441 4391 4487 4403
rect 4289 4359 4319 4362
rect 2949 4319 2961 4353
rect 3129 4319 3219 4353
rect 3387 4319 3477 4353
rect 3645 4319 3735 4353
rect 2949 4313 3777 4319
rect 2871 4310 2881 4313
rect 3763 4310 3777 4313
rect 3903 4313 3915 4359
rect 3981 4353 4319 4359
rect 4419 4359 4429 4362
rect 4556 4359 4644 5223
rect 4699 5179 4745 5191
rect 4699 4603 4705 5179
rect 4739 4603 4745 5179
rect 4684 4403 4694 4603
rect 4750 4403 4760 4603
rect 4699 4391 4745 4403
rect 4800 4359 4888 5223
rect 4957 5179 5003 5191
rect 4938 4979 4948 5179
rect 5012 4979 5022 5179
rect 4957 4403 4963 4979
rect 4997 4403 5003 4979
rect 4957 4391 5003 4403
rect 5065 4359 5153 5223
rect 5215 5179 5261 5191
rect 5215 4603 5221 5179
rect 5255 4603 5261 5179
rect 5200 4403 5210 4603
rect 5266 4403 5276 4603
rect 5215 4391 5261 4403
rect 5316 4362 5404 5223
rect 5473 5179 5519 5191
rect 5473 4827 5479 5179
rect 5513 4827 5519 5179
rect 5582 4830 5670 5223
rect 5731 5179 5777 5191
rect 5718 4979 5728 5179
rect 5780 4979 5790 5179
rect 5460 4727 5470 4827
rect 5522 4727 5532 4827
rect 5582 4730 5595 4830
rect 5647 4730 5670 4830
rect 5473 4403 5479 4727
rect 5513 4403 5519 4727
rect 5473 4391 5519 4403
rect 5316 4359 5326 4362
rect 3981 4319 3993 4353
rect 4161 4319 4251 4353
rect 3981 4313 4319 4319
rect 3903 4310 3913 4313
rect 4309 4310 4319 4313
rect 4419 4313 4431 4359
rect 4497 4353 5326 4359
rect 5451 4359 5461 4362
rect 5582 4359 5670 4730
rect 5731 4403 5737 4979
rect 5771 4403 5777 4979
rect 5731 4391 5777 4403
rect 5839 4833 5927 5223
rect 5839 4728 5857 4833
rect 5909 4728 5927 4833
rect 5989 5179 6035 5191
rect 5989 4827 5995 5179
rect 6029 4827 6035 5179
rect 5839 4362 5927 4728
rect 5976 4727 5986 4827
rect 6038 4727 6048 4827
rect 5989 4403 5995 4727
rect 6029 4403 6035 4727
rect 5989 4391 6035 4403
rect 5839 4359 5867 4362
rect 4497 4319 4509 4353
rect 4677 4319 4767 4353
rect 4935 4319 5025 4353
rect 5193 4319 5283 4353
rect 4497 4313 5326 4319
rect 4419 4310 4429 4313
rect 5320 4310 5326 4313
rect 5451 4313 5463 4359
rect 5529 4353 5867 4359
rect 5967 4359 5977 4362
rect 6113 4359 6201 5223
rect 6247 5179 6293 5191
rect 6247 4603 6253 5179
rect 6287 4603 6293 5179
rect 6232 4403 6242 4603
rect 6298 4403 6308 4603
rect 6247 4391 6293 4403
rect 6356 4362 6444 5223
rect 6505 5179 6551 5191
rect 6486 4979 6496 5179
rect 6560 4979 6570 5179
rect 6505 4403 6511 4979
rect 6545 4403 6551 4979
rect 6505 4391 6551 4403
rect 6356 4359 6383 4362
rect 5529 4319 5541 4353
rect 5709 4319 5799 4353
rect 5529 4313 5867 4319
rect 5451 4310 5461 4313
rect 5857 4310 5867 4313
rect 5967 4313 5979 4359
rect 6045 4353 6383 4359
rect 6483 4359 6493 4362
rect 6045 4319 6057 4353
rect 6225 4319 6315 4353
rect 6045 4313 6383 4319
rect 5967 4310 5977 4313
rect 6373 4310 6383 4313
rect 6483 4313 6495 4359
rect 6483 4310 6493 4313
rect 2206 4300 2251 4310
rect 94 4198 160 4210
rect 184 4084 755 4136
rect 855 4084 1529 4136
rect 1629 4084 2303 4136
rect 2403 4084 3077 4136
rect 3177 4084 3851 4136
rect 3951 4084 4625 4136
rect 4725 4084 5399 4136
rect 5499 4084 6173 4136
rect 6273 4084 6431 4136
rect 6531 4084 6541 4136
rect 184 2082 236 4084
rect 375 3939 497 3991
rect 597 3939 1271 3991
rect 1371 3939 2045 3991
rect 2145 3939 2819 3991
rect 2919 3939 3593 3991
rect 3693 3939 4367 3991
rect 4467 3939 5141 3991
rect 5241 3939 5915 3991
rect 6015 3939 6431 3991
rect 6531 3939 6541 3991
rect 439 3788 449 3791
rect 369 3782 449 3788
rect 549 3788 559 3791
rect 1371 3788 1381 3791
rect 369 3748 381 3782
rect 369 3742 449 3748
rect 426 3739 449 3742
rect 549 3742 561 3788
rect 627 3782 1381 3788
rect 1581 3788 1591 3791
rect 1987 3788 1997 3791
rect 627 3748 639 3782
rect 807 3748 897 3782
rect 1065 3748 1155 3782
rect 1323 3748 1381 3782
rect 627 3742 1381 3748
rect 549 3739 559 3742
rect 313 3698 359 3710
rect 313 3122 319 3698
rect 353 3122 359 3698
rect 426 3395 514 3739
rect 571 3698 617 3710
rect 571 3397 577 3698
rect 611 3397 617 3698
rect 426 3295 445 3395
rect 497 3295 514 3395
rect 558 3297 568 3397
rect 620 3297 630 3397
rect 300 2922 310 3122
rect 362 2922 372 3122
rect 313 2910 359 2922
rect 426 2878 514 3295
rect 571 2922 577 3297
rect 611 2922 617 3297
rect 571 2910 617 2922
rect 678 2878 766 3742
rect 829 3698 875 3710
rect 829 3123 835 3698
rect 869 3123 875 3698
rect 814 2923 824 3123
rect 880 2923 890 3123
rect 829 2922 835 2923
rect 869 2922 875 2923
rect 829 2910 875 2922
rect 927 2878 1015 3742
rect 1087 3698 1133 3710
rect 1068 3498 1078 3698
rect 1142 3498 1152 3698
rect 1087 2922 1093 3498
rect 1127 2922 1133 3498
rect 1087 2910 1133 2922
rect 1197 2878 1285 3742
rect 1371 3739 1381 3742
rect 1581 3742 1593 3788
rect 1659 3782 1997 3788
rect 2097 3788 2107 3791
rect 2935 3788 2945 3791
rect 1659 3748 1671 3782
rect 1839 3748 1929 3782
rect 1659 3742 1997 3748
rect 1581 3739 1591 3742
rect 1345 3698 1391 3710
rect 1345 3122 1351 3698
rect 1385 3122 1391 3698
rect 1330 2922 1340 3122
rect 1396 2922 1406 3122
rect 1345 2910 1391 2922
rect 1446 2878 1534 3739
rect 1603 3698 1649 3710
rect 1603 3397 1609 3698
rect 1643 3397 1649 3698
rect 1709 3398 1797 3742
rect 1963 3739 1997 3742
rect 2097 3742 2109 3788
rect 2175 3782 2945 3788
rect 3129 3788 3139 3791
rect 3535 3788 3545 3791
rect 2175 3748 2187 3782
rect 2355 3748 2445 3782
rect 2613 3748 2703 3782
rect 2871 3748 2945 3782
rect 2175 3742 2945 3748
rect 2097 3739 2107 3742
rect 1590 3297 1600 3397
rect 1652 3297 1662 3397
rect 1709 3298 1723 3398
rect 1775 3298 1797 3398
rect 1603 2922 1609 3297
rect 1643 2922 1649 3297
rect 1603 2910 1649 2922
rect 1709 2878 1797 3298
rect 1861 3698 1907 3710
rect 1861 3122 1867 3698
rect 1901 3122 1907 3698
rect 1963 3399 2051 3739
rect 1963 3299 1979 3399
rect 2031 3299 2051 3399
rect 2119 3698 2165 3710
rect 2119 3397 2125 3698
rect 2159 3397 2165 3698
rect 1848 2922 1858 3122
rect 1910 2922 1920 3122
rect 1861 2910 1907 2922
rect 1963 2878 2051 3299
rect 2106 3297 2116 3397
rect 2168 3297 2178 3397
rect 2119 2922 2125 3297
rect 2159 2922 2165 3297
rect 2119 2910 2165 2922
rect 2230 2878 2318 3742
rect 2377 3698 2423 3710
rect 2377 3122 2383 3698
rect 2417 3122 2423 3698
rect 2362 2922 2372 3122
rect 2428 2922 2438 3122
rect 2377 2910 2423 2922
rect 2483 2878 2571 3742
rect 2635 3698 2681 3710
rect 2616 3498 2626 3698
rect 2690 3498 2700 3698
rect 2635 2922 2641 3498
rect 2675 2922 2681 3498
rect 2635 2910 2681 2922
rect 2735 2878 2823 3742
rect 2935 3739 2945 3742
rect 3129 3742 3141 3788
rect 3207 3782 3545 3788
rect 3645 3788 3655 3791
rect 4483 3788 4493 3791
rect 3207 3748 3219 3782
rect 3387 3748 3477 3782
rect 3207 3742 3545 3748
rect 3129 3739 3139 3742
rect 2893 3698 2939 3710
rect 2893 3122 2899 3698
rect 2933 3122 2939 3698
rect 2878 2922 2888 3122
rect 2944 2922 2954 3122
rect 2893 2910 2939 2922
rect 3006 2878 3094 3739
rect 3151 3698 3197 3710
rect 3151 3397 3157 3698
rect 3191 3397 3197 3698
rect 3252 3397 3333 3742
rect 3512 3739 3545 3742
rect 3645 3742 3657 3788
rect 3723 3782 4493 3788
rect 4677 3788 4687 3791
rect 5083 3788 5093 3791
rect 3723 3748 3735 3782
rect 3903 3748 3993 3782
rect 4161 3748 4251 3782
rect 4419 3748 4493 3782
rect 3723 3742 4493 3748
rect 3645 3739 3655 3742
rect 3138 3297 3148 3397
rect 3200 3297 3210 3397
rect 3252 3297 3265 3397
rect 3317 3297 3333 3397
rect 3151 2922 3157 3297
rect 3191 2922 3197 3297
rect 3151 2910 3197 2922
rect 3252 2878 3333 3297
rect 3409 3698 3455 3710
rect 3409 3122 3415 3698
rect 3449 3122 3455 3698
rect 3512 3395 3593 3739
rect 3667 3698 3713 3710
rect 3667 3398 3673 3698
rect 3707 3398 3713 3698
rect 3512 3295 3527 3395
rect 3579 3295 3593 3395
rect 3654 3298 3664 3398
rect 3716 3298 3726 3398
rect 3396 2922 3406 3122
rect 3458 2922 3468 3122
rect 3409 2910 3455 2922
rect 3512 2878 3593 3295
rect 3667 2922 3673 3298
rect 3707 2922 3713 3298
rect 3667 2910 3713 2922
rect 3774 2878 3862 3742
rect 3925 3698 3971 3710
rect 3925 3122 3931 3698
rect 3965 3122 3971 3698
rect 3910 2922 3920 3122
rect 3976 2922 3986 3122
rect 3925 2910 3971 2922
rect 4030 2878 4118 3742
rect 4183 3698 4229 3710
rect 4164 3498 4174 3698
rect 4238 3498 4248 3698
rect 4183 2922 4189 3498
rect 4223 2922 4229 3498
rect 4183 2910 4229 2922
rect 4291 2878 4379 3742
rect 4483 3739 4493 3742
rect 4677 3742 4689 3788
rect 4755 3782 5093 3788
rect 5193 3788 5203 3791
rect 6031 3788 6041 3791
rect 4755 3748 4767 3782
rect 4935 3748 5025 3782
rect 4755 3742 5093 3748
rect 4677 3739 4687 3742
rect 4441 3698 4487 3710
rect 4441 3122 4447 3698
rect 4481 3122 4487 3698
rect 4426 2922 4436 3122
rect 4492 2922 4502 3122
rect 4441 2910 4487 2922
rect 4546 2878 4634 3739
rect 4699 3698 4745 3710
rect 4699 3397 4705 3698
rect 4739 3397 4745 3698
rect 4686 3297 4696 3397
rect 4748 3297 4758 3397
rect 4801 3395 4907 3742
rect 5056 3739 5093 3742
rect 5193 3742 5205 3788
rect 5271 3782 6041 3788
rect 6225 3788 6235 3791
rect 6373 3788 6383 3791
rect 5271 3748 5283 3782
rect 5451 3748 5541 3782
rect 5709 3748 5799 3782
rect 5967 3748 6041 3782
rect 5271 3742 6041 3748
rect 5193 3739 5203 3742
rect 4699 2922 4705 3297
rect 4739 2922 4745 3297
rect 4699 2910 4745 2922
rect 4801 3295 4823 3395
rect 4875 3295 4907 3395
rect 4801 2878 4907 3295
rect 4957 3698 5003 3710
rect 4957 3122 4963 3698
rect 4997 3122 5003 3698
rect 5056 3397 5162 3739
rect 5215 3698 5261 3710
rect 5215 3397 5221 3698
rect 5255 3397 5261 3698
rect 5056 3297 5078 3397
rect 5130 3297 5162 3397
rect 5202 3297 5212 3397
rect 5264 3297 5274 3397
rect 4944 2922 4954 3122
rect 5006 2922 5016 3122
rect 4957 2910 5003 2922
rect 5056 2878 5162 3297
rect 5215 2922 5221 3297
rect 5255 2922 5261 3297
rect 5215 2910 5261 2922
rect 5326 2878 5414 3742
rect 5473 3698 5519 3710
rect 5473 3122 5479 3698
rect 5513 3122 5519 3698
rect 5458 2922 5468 3122
rect 5524 2922 5534 3122
rect 5473 2910 5519 2922
rect 5582 2878 5670 3742
rect 5731 3698 5777 3710
rect 5712 3498 5722 3698
rect 5786 3498 5796 3698
rect 5731 2922 5737 3498
rect 5771 2922 5777 3498
rect 5731 2910 5777 2922
rect 5841 2878 5929 3742
rect 6031 3739 6041 3742
rect 6225 3742 6237 3788
rect 6303 3782 6383 3788
rect 6483 3788 6493 3791
rect 6303 3748 6315 3782
rect 6303 3742 6383 3748
rect 6225 3739 6235 3742
rect 6354 3739 6383 3742
rect 6483 3742 6495 3788
rect 6483 3739 6493 3742
rect 5989 3698 6035 3710
rect 5989 3122 5995 3698
rect 6029 3122 6035 3698
rect 5974 2922 5984 3122
rect 6040 2922 6050 3122
rect 5989 2910 6035 2922
rect 6101 2878 6189 3739
rect 6247 3698 6293 3710
rect 6247 3397 6253 3698
rect 6287 3397 6293 3698
rect 6354 3399 6442 3739
rect 6234 3297 6244 3397
rect 6296 3297 6306 3397
rect 6354 3299 6370 3399
rect 6422 3299 6442 3399
rect 6247 2922 6253 3297
rect 6287 2922 6293 3297
rect 6247 2910 6293 2922
rect 6354 2878 6442 3299
rect 6505 3698 6551 3710
rect 6505 3122 6511 3698
rect 6545 3122 6551 3698
rect 6492 2922 6502 3122
rect 6554 2922 6564 3122
rect 6505 2910 6551 2922
rect 369 2872 561 2878
rect 369 2838 381 2872
rect 549 2838 561 2872
rect 369 2832 561 2838
rect 627 2872 1593 2878
rect 627 2838 639 2872
rect 807 2838 897 2872
rect 1065 2838 1155 2872
rect 1323 2838 1413 2872
rect 1581 2838 1593 2872
rect 627 2832 1593 2838
rect 1659 2872 2109 2878
rect 1659 2838 1671 2872
rect 1839 2838 1929 2872
rect 2097 2838 2109 2872
rect 1659 2832 2109 2838
rect 2175 2872 3141 2878
rect 2175 2838 2187 2872
rect 2355 2838 2445 2872
rect 2613 2838 2703 2872
rect 2871 2838 2961 2872
rect 3129 2838 3141 2872
rect 2175 2832 3141 2838
rect 3207 2872 3657 2878
rect 3207 2838 3219 2872
rect 3387 2838 3477 2872
rect 3645 2838 3657 2872
rect 3207 2832 3657 2838
rect 3723 2872 4689 2878
rect 3723 2838 3735 2872
rect 3903 2838 3993 2872
rect 4161 2838 4251 2872
rect 4419 2838 4509 2872
rect 4677 2838 4689 2872
rect 3723 2832 4689 2838
rect 4755 2872 5205 2878
rect 4755 2838 4767 2872
rect 4935 2838 5025 2872
rect 5193 2838 5205 2872
rect 4755 2832 5205 2838
rect 5271 2872 6237 2878
rect 5271 2838 5283 2872
rect 5451 2838 5541 2872
rect 5709 2838 5799 2872
rect 5967 2838 6057 2872
rect 6225 2838 6237 2872
rect 5271 2832 6237 2838
rect 6303 2872 6495 2878
rect 6303 2838 6315 2872
rect 6483 2838 6495 2872
rect 6303 2832 6495 2838
rect 277 2663 6643 2669
rect 277 2551 290 2663
rect 6631 2551 6643 2663
rect 277 2545 6643 2551
rect 270 2502 821 2508
rect 270 2406 282 2502
rect 809 2406 821 2502
rect 270 2400 821 2406
rect 1177 2323 1297 2335
rect 184 2077 1028 2082
rect 184 2037 916 2077
rect 184 2030 449 2037
rect 418 2003 449 2030
rect 483 2003 549 2037
rect 583 2003 649 2037
rect 683 2003 749 2037
rect 783 2003 849 2037
rect 883 2003 916 2037
rect 418 1937 916 2003
rect 418 1903 449 1937
rect 483 1903 549 1937
rect 583 1903 649 1937
rect 683 1903 749 1937
rect 783 1903 849 1937
rect 883 1903 916 1937
rect 130 1890 262 1902
rect 126 1411 136 1890
rect 256 1411 266 1890
rect 418 1837 916 1903
rect 418 1803 449 1837
rect 483 1803 549 1837
rect 583 1803 649 1837
rect 683 1803 749 1837
rect 783 1803 849 1837
rect 883 1803 916 1837
rect 418 1737 916 1803
rect 418 1703 449 1737
rect 483 1703 549 1737
rect 583 1703 649 1737
rect 683 1703 749 1737
rect 783 1703 849 1737
rect 883 1703 916 1737
rect 418 1637 916 1703
rect 418 1603 449 1637
rect 483 1603 549 1637
rect 583 1603 649 1637
rect 683 1603 749 1637
rect 783 1603 849 1637
rect 883 1603 916 1637
rect 418 1537 916 1603
rect 418 1503 449 1537
rect 483 1503 549 1537
rect 583 1503 649 1537
rect 683 1503 749 1537
rect 783 1503 849 1537
rect 883 1503 916 1537
rect 418 1477 916 1503
rect 990 1477 1028 2077
rect 418 1472 1028 1477
rect 130 1399 262 1411
rect 221 1313 1070 1319
rect 221 1165 233 1313
rect 1058 1165 1070 1313
rect 1173 1280 1183 2323
rect 1291 1280 1301 2323
rect 2072 1922 7503 1928
rect 2072 1731 2084 1922
rect 7491 1731 7503 1922
rect 2072 1725 7503 1731
rect 2255 1646 3479 1652
rect 2255 1612 2267 1646
rect 2435 1612 2525 1646
rect 2693 1612 2783 1646
rect 2951 1612 3041 1646
rect 3209 1612 3299 1646
rect 3467 1612 3479 1646
rect 2255 1606 3479 1612
rect 3545 1646 4769 1652
rect 3545 1612 3557 1646
rect 3725 1612 3815 1646
rect 3983 1612 4073 1646
rect 4241 1612 4331 1646
rect 4499 1612 4589 1646
rect 4757 1612 4769 1646
rect 3545 1606 4769 1612
rect 4835 1646 6059 1652
rect 4835 1612 4847 1646
rect 5015 1612 5105 1646
rect 5273 1612 5363 1646
rect 5531 1612 5621 1646
rect 5789 1612 5879 1646
rect 6047 1612 6059 1646
rect 4835 1606 6059 1612
rect 6125 1646 7349 1652
rect 6125 1612 6137 1646
rect 6305 1612 6395 1646
rect 6563 1612 6653 1646
rect 6821 1612 6911 1646
rect 7079 1612 7169 1646
rect 7337 1612 7349 1646
rect 6125 1606 7349 1612
rect 2199 1562 2245 1574
rect 2186 1502 2196 1562
rect 2248 1502 2258 1562
rect 2199 1386 2205 1502
rect 2239 1386 2245 1502
rect 2199 1374 2245 1386
rect 2316 1342 2383 1606
rect 2457 1562 2503 1574
rect 2444 1502 2454 1562
rect 2506 1502 2516 1562
rect 2457 1386 2463 1502
rect 2497 1386 2503 1502
rect 2457 1374 2503 1386
rect 2574 1342 2641 1606
rect 2715 1562 2761 1606
rect 2715 1446 2721 1562
rect 2755 1446 2761 1562
rect 2702 1386 2712 1446
rect 2764 1386 2774 1446
rect 2702 1342 2774 1386
rect 2836 1342 2903 1606
rect 2973 1562 3019 1574
rect 2960 1502 2970 1562
rect 3022 1502 3032 1562
rect 2973 1386 2979 1502
rect 3013 1386 3019 1502
rect 2973 1374 3019 1386
rect 3093 1342 3160 1606
rect 3231 1562 3277 1606
rect 3231 1446 3237 1562
rect 3271 1446 3277 1562
rect 3218 1386 3228 1446
rect 3280 1386 3290 1446
rect 3218 1342 3290 1386
rect 3353 1342 3420 1606
rect 3489 1562 3535 1574
rect 3476 1502 3486 1562
rect 3538 1502 3548 1562
rect 3489 1386 3495 1502
rect 3529 1386 3535 1502
rect 3489 1374 3535 1386
rect 3605 1342 3672 1606
rect 3747 1562 3793 1574
rect 3734 1502 3744 1562
rect 3796 1502 3806 1562
rect 3747 1386 3753 1502
rect 3787 1386 3793 1502
rect 3747 1374 3793 1386
rect 3859 1342 3926 1606
rect 4005 1562 4051 1606
rect 4005 1446 4011 1562
rect 4045 1446 4051 1562
rect 3992 1386 4002 1446
rect 4054 1386 4064 1446
rect 3992 1342 4064 1386
rect 4120 1342 4187 1606
rect 4263 1562 4309 1574
rect 4250 1502 4260 1562
rect 4312 1502 4322 1562
rect 4263 1386 4269 1502
rect 4303 1386 4309 1502
rect 4263 1374 4309 1386
rect 4373 1342 4440 1606
rect 4521 1562 4567 1606
rect 4521 1446 4527 1562
rect 4561 1446 4567 1562
rect 4508 1386 4518 1446
rect 4570 1386 4580 1446
rect 4508 1342 4580 1386
rect 4635 1342 4702 1606
rect 4779 1562 4825 1574
rect 4766 1502 4776 1562
rect 4828 1502 4838 1562
rect 4779 1386 4785 1502
rect 4819 1386 4825 1502
rect 4779 1374 4825 1386
rect 4893 1342 4960 1606
rect 5037 1562 5083 1574
rect 5024 1502 5034 1562
rect 5086 1502 5096 1562
rect 5037 1386 5043 1502
rect 5077 1386 5083 1502
rect 5037 1374 5083 1386
rect 5150 1342 5217 1606
rect 5295 1562 5341 1606
rect 5295 1446 5301 1562
rect 5335 1446 5341 1562
rect 5282 1386 5292 1446
rect 5344 1386 5354 1446
rect 5282 1342 5354 1386
rect 5411 1342 5478 1606
rect 5553 1562 5599 1574
rect 5540 1502 5550 1562
rect 5602 1502 5612 1562
rect 5553 1386 5559 1502
rect 5593 1386 5599 1502
rect 5553 1374 5599 1386
rect 5670 1342 5737 1606
rect 5811 1562 5857 1606
rect 5811 1446 5817 1562
rect 5851 1446 5857 1562
rect 5798 1386 5808 1446
rect 5860 1386 5870 1446
rect 5798 1342 5870 1386
rect 5920 1342 5987 1606
rect 6069 1562 6115 1574
rect 6056 1502 6066 1562
rect 6118 1502 6128 1562
rect 6069 1386 6075 1502
rect 6109 1386 6115 1502
rect 6069 1374 6115 1386
rect 6180 1342 6247 1606
rect 6327 1562 6373 1574
rect 6314 1502 6324 1562
rect 6376 1502 6386 1562
rect 6327 1386 6333 1502
rect 6367 1386 6373 1502
rect 6327 1374 6373 1386
rect 6442 1342 6509 1606
rect 6585 1562 6631 1606
rect 6585 1446 6591 1562
rect 6625 1446 6631 1562
rect 6572 1386 6582 1446
rect 6634 1386 6644 1446
rect 6572 1342 6644 1386
rect 6702 1342 6769 1606
rect 6843 1562 6889 1574
rect 6830 1502 6840 1562
rect 6892 1502 6902 1562
rect 6843 1386 6849 1502
rect 6883 1386 6889 1502
rect 6843 1374 6889 1386
rect 6961 1342 7028 1606
rect 7101 1562 7147 1606
rect 7101 1446 7107 1562
rect 7141 1446 7147 1562
rect 7088 1386 7098 1446
rect 7150 1386 7160 1446
rect 7088 1342 7160 1386
rect 7228 1342 7295 1606
rect 7359 1562 7405 1574
rect 7346 1502 7356 1562
rect 7408 1502 7418 1562
rect 7359 1446 7365 1502
rect 7399 1446 7405 1502
rect 7346 1386 7356 1446
rect 7408 1386 7418 1446
rect 7359 1374 7405 1386
rect 2255 1336 3479 1342
rect 2255 1302 2267 1336
rect 2435 1302 2525 1336
rect 2693 1302 2783 1336
rect 2951 1302 3041 1336
rect 3209 1302 3299 1336
rect 3467 1302 3479 1336
rect 2255 1296 3479 1302
rect 3545 1336 4769 1342
rect 3545 1302 3557 1336
rect 3725 1302 3815 1336
rect 3983 1302 4073 1336
rect 4241 1302 4331 1336
rect 4499 1302 4589 1336
rect 4757 1302 4769 1336
rect 3545 1296 4769 1302
rect 4835 1336 6059 1342
rect 4835 1302 4847 1336
rect 5015 1302 5105 1336
rect 5273 1302 5363 1336
rect 5531 1302 5621 1336
rect 5789 1302 5879 1336
rect 6047 1302 6059 1336
rect 4835 1296 6059 1302
rect 6125 1336 7349 1342
rect 6125 1302 6137 1336
rect 6305 1302 6395 1336
rect 6563 1302 6653 1336
rect 6821 1302 6911 1336
rect 7079 1302 7169 1336
rect 7337 1302 7349 1336
rect 6125 1296 7349 1302
rect 1177 1268 1297 1280
rect 221 1159 1070 1165
rect 260 873 270 894
rect 195 867 270 873
rect 629 873 639 894
rect 714 873 724 894
rect 629 867 724 873
rect 1083 873 1093 894
rect 1753 873 7419 874
rect 1083 868 7419 873
rect 1083 867 2583 868
rect 195 833 263 867
rect 631 833 721 867
rect 1089 833 1388 867
rect 1556 833 1646 867
rect 1814 834 2583 867
rect 2951 834 3873 868
rect 4241 834 5163 868
rect 5531 834 6453 868
rect 6821 834 7034 868
rect 7402 834 7419 868
rect 1814 833 7419 834
rect 195 829 270 833
rect 629 829 724 833
rect 1083 829 7419 833
rect 195 828 7419 829
rect 195 827 2401 828
rect 195 774 241 827
rect 195 698 201 774
rect 235 698 241 774
rect 195 686 241 698
rect 310 645 592 827
rect 653 774 699 786
rect 640 698 650 774
rect 702 698 712 774
rect 653 686 699 698
rect 757 645 1039 827
rect 1111 774 1157 827
rect 1320 774 1366 786
rect 1111 698 1117 774
rect 1151 698 1157 774
rect 1111 686 1157 698
rect 251 639 643 645
rect 251 605 263 639
rect 631 605 643 639
rect 251 599 643 605
rect 709 639 1101 645
rect 709 605 721 639
rect 1089 605 1101 639
rect 1301 634 1311 774
rect 1375 634 1385 774
rect 709 599 1101 605
rect 1320 598 1326 634
rect 1360 598 1366 634
rect 1320 586 1366 598
rect 1419 545 1537 827
rect 1578 774 1624 786
rect 1578 738 1584 774
rect 1618 738 1624 774
rect 1565 598 1575 738
rect 1627 598 1637 738
rect 1578 586 1624 598
rect 1671 545 1789 827
rect 1836 774 1882 786
rect 2515 775 2561 787
rect 1817 634 1827 774
rect 1891 634 1901 774
rect 2515 722 2521 775
rect 2555 722 2561 775
rect 1836 598 1842 634
rect 1876 598 1882 634
rect 2502 599 2512 722
rect 2564 599 2574 722
rect 1836 586 1882 598
rect 2515 587 2561 599
rect 2621 546 2900 828
rect 2973 775 3019 787
rect 3805 775 3851 787
rect 2960 662 2970 775
rect 3022 662 3032 775
rect 3805 722 3811 775
rect 3845 722 3851 775
rect 2973 599 2979 662
rect 3013 599 3019 662
rect 3792 599 3802 722
rect 3854 599 3864 722
rect 2973 587 3019 599
rect 3805 587 3851 599
rect 3919 546 4198 828
rect 4263 775 4309 787
rect 5095 775 5141 787
rect 4250 662 4260 775
rect 4312 662 4322 775
rect 5095 722 5101 775
rect 5135 722 5141 775
rect 4263 599 4269 662
rect 4303 599 4309 662
rect 5082 599 5092 722
rect 5144 599 5154 722
rect 4263 587 4309 599
rect 5095 587 5141 599
rect 5200 546 5479 828
rect 5553 775 5599 787
rect 6385 775 6431 787
rect 5540 662 5550 775
rect 5602 662 5612 775
rect 6385 723 6391 775
rect 6425 723 6431 775
rect 5553 599 5559 662
rect 5593 599 5599 662
rect 6372 599 6382 723
rect 6434 599 6444 723
rect 5553 587 5599 599
rect 6385 587 6431 599
rect 6510 546 6789 828
rect 6843 775 6889 787
rect 6966 775 7012 787
rect 6830 652 6840 775
rect 6892 652 6902 775
rect 6966 722 6972 775
rect 7006 722 7012 775
rect 6843 599 6849 652
rect 6883 599 6889 652
rect 6953 599 6963 722
rect 7015 599 7025 722
rect 6843 587 6889 599
rect 6966 587 7012 599
rect 7086 546 7365 828
rect 7424 775 7470 787
rect 7411 652 7421 775
rect 7473 652 7483 775
rect 7424 599 7430 652
rect 7464 599 7470 652
rect 7424 587 7470 599
rect 1376 539 1568 545
rect 1376 505 1388 539
rect 1556 505 1568 539
rect 1376 499 1568 505
rect 1634 539 1826 545
rect 1634 505 1646 539
rect 1814 505 1826 539
rect 1634 499 1826 505
rect 2571 540 2963 546
rect 2571 506 2583 540
rect 2951 506 2963 540
rect 2571 500 2963 506
rect 3861 540 4253 546
rect 3861 506 3873 540
rect 4241 506 4253 540
rect 3861 500 4253 506
rect 5151 540 5543 546
rect 5151 506 5163 540
rect 5531 506 5543 540
rect 5151 500 5543 506
rect 6441 540 6833 546
rect 6441 506 6453 540
rect 6821 506 6833 540
rect 6441 500 6833 506
rect 7022 540 7414 546
rect 7022 506 7034 540
rect 7402 506 7414 540
rect 7022 500 7414 506
rect 1005 445 2015 447
rect 12 441 2015 445
rect 12 439 1017 441
rect 12 307 24 439
rect 12 306 1017 307
rect 2003 306 2015 441
rect 6194 334 6252 338
rect 12 301 2015 306
rect 1005 300 2015 301
rect 2502 328 6167 334
rect 13 228 2016 234
rect 13 80 25 228
rect 2004 80 2016 228
rect 2502 189 2514 328
rect 2502 183 6167 189
rect 7521 183 7531 334
rect 6194 179 6252 183
rect 13 74 2016 80
<< via1 >>
rect 97 5430 6675 5604
rect 100 5196 154 5348
rect 304 4979 319 5179
rect 319 4979 353 5179
rect 353 4979 368 5179
rect 566 4403 577 4603
rect 577 4403 611 4603
rect 611 4403 622 4603
rect 1084 4979 1093 5179
rect 1093 4979 1127 5179
rect 1127 4979 1136 5179
rect 826 4727 835 4827
rect 835 4727 869 4827
rect 869 4727 878 4827
rect 950 4727 1002 4827
rect 100 4210 154 4358
rect 707 4353 807 4362
rect 1215 4727 1267 4827
rect 1342 4727 1351 4827
rect 1351 4727 1385 4827
rect 1385 4727 1394 4827
rect 707 4319 807 4353
rect 707 4310 807 4319
rect 1223 4353 1323 4362
rect 1598 4403 1609 4603
rect 1609 4403 1643 4603
rect 1643 4403 1654 4603
rect 1852 4979 1867 5179
rect 1867 4979 1901 5179
rect 1901 4979 1916 5179
rect 2114 4403 2125 4603
rect 2125 4403 2159 4603
rect 2159 4403 2170 4603
rect 2632 4979 2641 5179
rect 2641 4979 2675 5179
rect 2675 4979 2684 5179
rect 2374 4727 2383 4827
rect 2383 4727 2417 4827
rect 2417 4727 2426 4827
rect 2497 4728 2549 4828
rect 1223 4319 1323 4353
rect 1223 4310 1323 4319
rect 2229 4353 2355 4362
rect 2759 4726 2811 4826
rect 2890 4727 2899 4827
rect 2899 4727 2933 4827
rect 2933 4727 2942 4827
rect 2229 4319 2355 4353
rect 2229 4310 2355 4319
rect 2771 4353 2871 4362
rect 3146 4403 3157 4603
rect 3157 4403 3191 4603
rect 3191 4403 3202 4603
rect 3400 4979 3415 5179
rect 3415 4979 3449 5179
rect 3449 4979 3464 5179
rect 3662 4403 3673 4603
rect 3673 4403 3707 4603
rect 3707 4403 3718 4603
rect 3922 4727 3931 4827
rect 3931 4727 3965 4827
rect 3965 4727 3974 4827
rect 4179 4979 4189 5179
rect 4189 4979 4223 5179
rect 4223 4979 4231 5179
rect 4052 4725 4104 4825
rect 2771 4319 2871 4353
rect 2771 4310 2871 4319
rect 3777 4353 3903 4362
rect 4304 4728 4356 4828
rect 4438 4727 4447 4827
rect 4447 4727 4481 4827
rect 4481 4727 4490 4827
rect 3777 4319 3903 4353
rect 3777 4310 3903 4319
rect 4319 4353 4419 4362
rect 4694 4403 4705 4603
rect 4705 4403 4739 4603
rect 4739 4403 4750 4603
rect 4948 4979 4963 5179
rect 4963 4979 4997 5179
rect 4997 4979 5012 5179
rect 5210 4403 5221 4603
rect 5221 4403 5255 4603
rect 5255 4403 5266 4603
rect 5728 4979 5737 5179
rect 5737 4979 5771 5179
rect 5771 4979 5780 5179
rect 5470 4727 5479 4827
rect 5479 4727 5513 4827
rect 5513 4727 5522 4827
rect 5595 4730 5647 4830
rect 4319 4319 4419 4353
rect 4319 4310 4419 4319
rect 5326 4353 5451 4362
rect 5857 4728 5909 4833
rect 5986 4727 5995 4827
rect 5995 4727 6029 4827
rect 6029 4727 6038 4827
rect 5326 4319 5451 4353
rect 5326 4310 5451 4319
rect 5867 4353 5967 4362
rect 6242 4403 6253 4603
rect 6253 4403 6287 4603
rect 6287 4403 6298 4603
rect 6496 4979 6511 5179
rect 6511 4979 6545 5179
rect 6545 4979 6560 5179
rect 5867 4319 5967 4353
rect 5867 4310 5967 4319
rect 6383 4353 6483 4362
rect 6383 4319 6483 4353
rect 6383 4310 6483 4319
rect 755 4084 855 4136
rect 1529 4084 1629 4136
rect 2303 4084 2403 4136
rect 3077 4084 3177 4136
rect 3851 4084 3951 4136
rect 4625 4084 4725 4136
rect 5399 4084 5499 4136
rect 6173 4084 6273 4136
rect 6431 4084 6531 4136
rect 497 3939 597 3991
rect 1271 3939 1371 3991
rect 2045 3939 2145 3991
rect 2819 3939 2919 3991
rect 3593 3939 3693 3991
rect 4367 3939 4467 3991
rect 5141 3939 5241 3991
rect 5915 3939 6015 3991
rect 6431 3939 6531 3991
rect 449 3782 549 3791
rect 449 3748 549 3782
rect 449 3739 549 3748
rect 1381 3782 1581 3791
rect 1381 3748 1413 3782
rect 1413 3748 1581 3782
rect 445 3295 497 3395
rect 568 3297 577 3397
rect 577 3297 611 3397
rect 611 3297 620 3397
rect 310 2922 319 3122
rect 319 2922 353 3122
rect 353 2922 362 3122
rect 824 2923 835 3123
rect 835 2923 869 3123
rect 869 2923 880 3123
rect 1078 3498 1093 3698
rect 1093 3498 1127 3698
rect 1127 3498 1142 3698
rect 1381 3739 1581 3748
rect 1997 3782 2097 3791
rect 1997 3748 2097 3782
rect 1340 2922 1351 3122
rect 1351 2922 1385 3122
rect 1385 2922 1396 3122
rect 1997 3739 2097 3748
rect 2945 3782 3129 3791
rect 2945 3748 2961 3782
rect 2961 3748 3129 3782
rect 1600 3297 1609 3397
rect 1609 3297 1643 3397
rect 1643 3297 1652 3397
rect 1723 3298 1775 3398
rect 1979 3299 2031 3399
rect 1858 2922 1867 3122
rect 1867 2922 1901 3122
rect 1901 2922 1910 3122
rect 2116 3297 2125 3397
rect 2125 3297 2159 3397
rect 2159 3297 2168 3397
rect 2372 2922 2383 3122
rect 2383 2922 2417 3122
rect 2417 2922 2428 3122
rect 2626 3498 2641 3698
rect 2641 3498 2675 3698
rect 2675 3498 2690 3698
rect 2945 3739 3129 3748
rect 3545 3782 3645 3791
rect 3545 3748 3645 3782
rect 2888 2922 2899 3122
rect 2899 2922 2933 3122
rect 2933 2922 2944 3122
rect 3545 3739 3645 3748
rect 4493 3782 4677 3791
rect 4493 3748 4509 3782
rect 4509 3748 4677 3782
rect 3148 3297 3157 3397
rect 3157 3297 3191 3397
rect 3191 3297 3200 3397
rect 3265 3297 3317 3397
rect 3527 3295 3579 3395
rect 3664 3298 3673 3398
rect 3673 3298 3707 3398
rect 3707 3298 3716 3398
rect 3406 2922 3415 3122
rect 3415 2922 3449 3122
rect 3449 2922 3458 3122
rect 3920 2922 3931 3122
rect 3931 2922 3965 3122
rect 3965 2922 3976 3122
rect 4174 3498 4189 3698
rect 4189 3498 4223 3698
rect 4223 3498 4238 3698
rect 4493 3739 4677 3748
rect 5093 3782 5193 3791
rect 5093 3748 5193 3782
rect 4436 2922 4447 3122
rect 4447 2922 4481 3122
rect 4481 2922 4492 3122
rect 4696 3297 4705 3397
rect 4705 3297 4739 3397
rect 4739 3297 4748 3397
rect 5093 3739 5193 3748
rect 6041 3782 6225 3791
rect 6041 3748 6057 3782
rect 6057 3748 6225 3782
rect 4823 3295 4875 3395
rect 5078 3297 5130 3397
rect 5212 3297 5221 3397
rect 5221 3297 5255 3397
rect 5255 3297 5264 3397
rect 4954 2922 4963 3122
rect 4963 2922 4997 3122
rect 4997 2922 5006 3122
rect 5468 2922 5479 3122
rect 5479 2922 5513 3122
rect 5513 2922 5524 3122
rect 5722 3498 5737 3698
rect 5737 3498 5771 3698
rect 5771 3498 5786 3698
rect 6041 3739 6225 3748
rect 6383 3782 6483 3791
rect 6383 3748 6483 3782
rect 6383 3739 6483 3748
rect 5984 2922 5995 3122
rect 5995 2922 6029 3122
rect 6029 2922 6040 3122
rect 6244 3297 6253 3397
rect 6253 3297 6287 3397
rect 6287 3297 6296 3397
rect 6370 3299 6422 3399
rect 6502 2922 6511 3122
rect 6511 2922 6545 3122
rect 6545 2922 6554 3122
rect 290 2551 6631 2663
rect 282 2406 809 2502
rect 916 2037 990 2077
rect 916 2003 949 2037
rect 949 2003 983 2037
rect 983 2003 990 2037
rect 916 1937 990 2003
rect 916 1903 949 1937
rect 949 1903 983 1937
rect 983 1903 990 1937
rect 136 1411 256 1890
rect 916 1837 990 1903
rect 916 1803 949 1837
rect 949 1803 983 1837
rect 983 1803 990 1837
rect 916 1737 990 1803
rect 916 1703 949 1737
rect 949 1703 983 1737
rect 983 1703 990 1737
rect 916 1637 990 1703
rect 916 1603 949 1637
rect 949 1603 983 1637
rect 983 1603 990 1637
rect 916 1537 990 1603
rect 916 1503 949 1537
rect 949 1503 983 1537
rect 983 1503 990 1537
rect 916 1477 990 1503
rect 233 1165 1058 1313
rect 1183 1280 1291 2323
rect 2084 1731 7491 1922
rect 2196 1502 2205 1562
rect 2205 1502 2239 1562
rect 2239 1502 2248 1562
rect 2454 1502 2463 1562
rect 2463 1502 2497 1562
rect 2497 1502 2506 1562
rect 2712 1386 2721 1446
rect 2721 1386 2755 1446
rect 2755 1386 2764 1446
rect 2970 1502 2979 1562
rect 2979 1502 3013 1562
rect 3013 1502 3022 1562
rect 3228 1386 3237 1446
rect 3237 1386 3271 1446
rect 3271 1386 3280 1446
rect 3486 1502 3495 1562
rect 3495 1502 3529 1562
rect 3529 1502 3538 1562
rect 3744 1502 3753 1562
rect 3753 1502 3787 1562
rect 3787 1502 3796 1562
rect 4002 1386 4011 1446
rect 4011 1386 4045 1446
rect 4045 1386 4054 1446
rect 4260 1502 4269 1562
rect 4269 1502 4303 1562
rect 4303 1502 4312 1562
rect 4518 1386 4527 1446
rect 4527 1386 4561 1446
rect 4561 1386 4570 1446
rect 4776 1502 4785 1562
rect 4785 1502 4819 1562
rect 4819 1502 4828 1562
rect 5034 1502 5043 1562
rect 5043 1502 5077 1562
rect 5077 1502 5086 1562
rect 5292 1386 5301 1446
rect 5301 1386 5335 1446
rect 5335 1386 5344 1446
rect 5550 1502 5559 1562
rect 5559 1502 5593 1562
rect 5593 1502 5602 1562
rect 5808 1386 5817 1446
rect 5817 1386 5851 1446
rect 5851 1386 5860 1446
rect 6066 1502 6075 1562
rect 6075 1502 6109 1562
rect 6109 1502 6118 1562
rect 6324 1502 6333 1562
rect 6333 1502 6367 1562
rect 6367 1502 6376 1562
rect 6582 1386 6591 1446
rect 6591 1386 6625 1446
rect 6625 1386 6634 1446
rect 6840 1502 6849 1562
rect 6849 1502 6883 1562
rect 6883 1502 6892 1562
rect 7098 1386 7107 1446
rect 7107 1386 7141 1446
rect 7141 1386 7150 1446
rect 7356 1502 7365 1562
rect 7365 1502 7399 1562
rect 7399 1502 7408 1562
rect 7356 1386 7365 1446
rect 7365 1386 7399 1446
rect 7399 1386 7408 1446
rect 270 867 629 894
rect 724 867 1083 894
rect 270 833 629 867
rect 724 833 1083 867
rect 270 829 629 833
rect 724 829 1083 833
rect 650 698 659 774
rect 659 698 693 774
rect 693 698 702 774
rect 1311 634 1326 774
rect 1326 634 1360 774
rect 1360 634 1375 774
rect 1575 598 1584 738
rect 1584 598 1618 738
rect 1618 598 1627 738
rect 1827 634 1842 774
rect 1842 634 1876 774
rect 1876 634 1891 774
rect 2512 599 2521 722
rect 2521 599 2555 722
rect 2555 599 2564 722
rect 2970 662 2979 775
rect 2979 662 3013 775
rect 3013 662 3022 775
rect 3802 599 3811 722
rect 3811 599 3845 722
rect 3845 599 3854 722
rect 4260 662 4269 775
rect 4269 662 4303 775
rect 4303 662 4312 775
rect 5092 599 5101 722
rect 5101 599 5135 722
rect 5135 599 5144 722
rect 5550 662 5559 775
rect 5559 662 5593 775
rect 5593 662 5602 775
rect 6382 599 6391 723
rect 6391 599 6425 723
rect 6425 599 6434 723
rect 6840 652 6849 775
rect 6849 652 6883 775
rect 6883 652 6892 775
rect 6963 599 6972 722
rect 6972 599 7006 722
rect 7006 599 7015 722
rect 7421 652 7430 775
rect 7430 652 7464 775
rect 7464 652 7473 775
rect 1017 439 1916 441
rect 24 406 1916 439
rect 1916 406 2003 441
rect 24 307 2003 406
rect 1017 306 2003 307
rect 6167 328 7521 334
rect 25 80 2004 228
rect 2514 189 7509 328
rect 7509 189 7521 328
rect 6167 183 7521 189
<< metal2 >>
rect -52 5604 6675 5614
rect -52 5430 97 5604
rect -52 5420 6675 5430
rect 100 5348 154 5420
rect 100 4358 154 5196
rect 304 5179 368 5189
rect 304 4969 368 4979
rect 1084 5179 1136 5420
rect 1084 4969 1136 4979
rect 1852 5179 1916 5189
rect 1852 4969 1916 4979
rect 2632 5179 2684 5420
rect 2632 4969 2684 4979
rect 3400 5179 3464 5189
rect 3400 4969 3464 4979
rect 4179 5179 4231 5420
rect 4179 4969 4231 4979
rect 4948 5179 5012 5189
rect 4948 4969 5012 4979
rect 5728 5179 5780 5420
rect 5728 4969 5780 4979
rect 6496 5179 6560 5189
rect 6496 4969 6560 4979
rect 2497 4837 2549 4838
rect 4304 4837 4356 4838
rect 5595 4837 5647 4840
rect 5857 4837 5909 4838
rect 826 4833 6834 4837
rect 826 4830 5857 4833
rect 826 4828 5595 4830
rect 826 4827 2497 4828
rect 878 4727 950 4827
rect 1002 4727 1215 4827
rect 1267 4727 1342 4827
rect 1394 4727 2374 4827
rect 2426 4728 2497 4827
rect 2549 4827 4304 4828
rect 2549 4826 2890 4827
rect 2549 4728 2759 4826
rect 2426 4727 2759 4728
rect 826 4726 2759 4727
rect 2811 4727 2890 4826
rect 2942 4727 3922 4827
rect 3974 4825 4304 4827
rect 3974 4727 4052 4825
rect 2811 4726 4052 4727
rect 826 4725 4052 4726
rect 4104 4728 4304 4825
rect 4356 4827 5595 4828
rect 4356 4728 4438 4827
rect 4104 4727 4438 4728
rect 4490 4727 5470 4827
rect 5522 4730 5595 4827
rect 5647 4730 5857 4830
rect 5522 4728 5857 4730
rect 5909 4827 6834 4833
rect 5909 4728 5986 4827
rect 5522 4727 5986 4728
rect 6038 4727 6834 4827
rect 4104 4725 6834 4727
rect 826 4717 6834 4725
rect 2759 4716 2811 4717
rect 4052 4715 4104 4717
rect 566 4603 622 4613
rect 566 4393 622 4403
rect 1598 4603 1654 4613
rect 1598 4393 1654 4403
rect 2114 4603 2170 4613
rect 2114 4393 2170 4403
rect 3146 4603 3202 4613
rect 3146 4393 3202 4403
rect 3662 4603 3718 4613
rect 3662 4393 3718 4403
rect 4694 4603 4750 4613
rect 4694 4393 4750 4403
rect 5210 4603 5266 4613
rect 5210 4393 5266 4403
rect 6242 4603 6298 4613
rect 6242 4393 6298 4403
rect 707 4362 807 4372
rect 707 4300 807 4310
rect 1223 4362 1323 4372
rect 1223 4300 1323 4310
rect 2223 4362 2355 4372
rect 2223 4310 2229 4362
rect 2223 4300 2355 4310
rect 2771 4362 2871 4372
rect 2771 4300 2871 4310
rect 3777 4362 3903 4372
rect 3777 4300 3903 4310
rect 4319 4362 4419 4372
rect 4319 4300 4419 4310
rect 5326 4362 5451 4372
rect 5326 4300 5451 4310
rect 5867 4362 5967 4372
rect 5867 4300 5967 4310
rect 6383 4362 6483 4372
rect 6383 4300 6483 4310
rect 100 2673 154 4210
rect 755 4146 807 4300
rect 755 4136 855 4146
rect 755 4074 855 4084
rect 1271 4001 1323 4300
rect 2303 4146 2355 4300
rect 1529 4136 1629 4146
rect 1529 4074 1629 4084
rect 2303 4136 2403 4146
rect 2303 4074 2403 4084
rect 497 3991 597 4001
rect 497 3929 597 3939
rect 1271 3991 1371 4001
rect 1271 3929 1371 3939
rect 497 3801 549 3929
rect 1529 3801 1581 4074
rect 2819 4001 2871 4300
rect 3851 4146 3903 4300
rect 3077 4136 3177 4146
rect 3077 4074 3177 4084
rect 3851 4136 3951 4146
rect 3851 4074 3951 4084
rect 2045 3991 2145 4001
rect 2045 3929 2145 3939
rect 2819 3991 2919 4001
rect 2819 3929 2919 3939
rect 2045 3801 2097 3929
rect 3077 3801 3129 4074
rect 4367 4001 4419 4300
rect 5399 4146 5451 4300
rect 4625 4136 4725 4146
rect 4625 4074 4725 4084
rect 5399 4136 5499 4146
rect 5399 4074 5499 4084
rect 3593 3991 3693 4001
rect 3593 3929 3693 3939
rect 4367 3991 4467 4001
rect 4367 3929 4467 3939
rect 3593 3801 3645 3929
rect 4625 3801 4677 4074
rect 5915 4001 5967 4300
rect 6431 4146 6483 4300
rect 6173 4136 6273 4146
rect 6173 4074 6273 4084
rect 6431 4136 6531 4146
rect 6431 4074 6531 4084
rect 5141 3991 5241 4001
rect 5141 3929 5241 3939
rect 5915 3991 6015 4001
rect 5915 3929 6015 3939
rect 5141 3801 5193 3929
rect 6173 3801 6225 4074
rect 6431 3991 6531 4001
rect 6431 3929 6531 3939
rect 6431 3801 6483 3929
rect 449 3791 549 3801
rect 449 3729 549 3739
rect 1381 3791 1581 3801
rect 1381 3729 1581 3739
rect 1997 3791 2097 3801
rect 1997 3729 2097 3739
rect 2945 3791 3129 3801
rect 2945 3729 3129 3739
rect 3545 3791 3645 3801
rect 3545 3729 3645 3739
rect 4493 3791 4677 3801
rect 4493 3729 4677 3739
rect 5093 3791 5193 3801
rect 5093 3729 5193 3739
rect 6041 3791 6225 3801
rect 6041 3729 6225 3739
rect 6383 3791 6483 3801
rect 6383 3729 6483 3739
rect 1078 3698 1142 3708
rect 1078 3488 1142 3498
rect 2626 3698 2690 3708
rect 2626 3488 2690 3498
rect 4174 3698 4238 3708
rect 4174 3488 4238 3498
rect 5722 3698 5786 3708
rect 5722 3488 5786 3498
rect 1723 3407 1775 3408
rect 1979 3407 2031 3409
rect 3664 3407 3716 3408
rect 6370 3407 6422 3409
rect 6714 3407 6834 4717
rect 421 3399 6834 3407
rect 421 3398 1979 3399
rect 421 3397 1723 3398
rect 421 3395 568 3397
rect 421 3295 445 3395
rect 497 3297 568 3395
rect 620 3297 1600 3397
rect 1652 3298 1723 3397
rect 1775 3299 1979 3398
rect 2031 3398 6370 3399
rect 2031 3397 3664 3398
rect 2031 3299 2116 3397
rect 1775 3298 2116 3299
rect 1652 3297 2116 3298
rect 2168 3297 3148 3397
rect 3200 3297 3265 3397
rect 3317 3395 3664 3397
rect 3317 3297 3527 3395
rect 497 3295 3527 3297
rect 3579 3298 3664 3395
rect 3716 3397 6370 3398
rect 3716 3298 4696 3397
rect 3579 3297 4696 3298
rect 4748 3395 5078 3397
rect 4748 3297 4823 3395
rect 3579 3295 4823 3297
rect 4875 3297 5078 3395
rect 5130 3297 5212 3397
rect 5264 3297 6244 3397
rect 6296 3299 6370 3397
rect 6422 3299 6834 3399
rect 6296 3297 6834 3299
rect 4875 3295 6834 3297
rect 421 3287 6834 3295
rect 445 3285 497 3287
rect 3527 3285 3579 3287
rect 4823 3285 4875 3287
rect 310 3122 362 3132
rect 310 2673 362 2922
rect 824 3123 880 3133
rect 824 2913 880 2923
rect 1340 3122 1396 3132
rect 1340 2912 1396 2922
rect 1858 3122 1910 3132
rect 1858 2673 1910 2922
rect 2372 3122 2428 3132
rect 2372 2912 2428 2922
rect 2888 3122 2944 3132
rect 2888 2912 2944 2922
rect 3406 3122 3458 3132
rect 3406 2673 3458 2922
rect 3920 3122 3976 3132
rect 3920 2912 3976 2922
rect 4436 3122 4492 3132
rect 4436 2912 4492 2922
rect 4954 3122 5006 3132
rect 4954 2673 5006 2922
rect 5468 3122 5524 3132
rect 5468 2912 5524 2922
rect 5984 3122 6040 3132
rect 5984 2912 6040 2922
rect 6502 3122 6554 3132
rect 6502 2673 6554 2922
rect 100 2663 6631 2673
rect 100 2619 290 2663
rect 277 2551 290 2619
rect 277 2541 6631 2551
rect 277 2502 809 2541
rect 277 2406 282 2502
rect 277 2396 809 2406
rect 1161 2323 1315 2541
rect 916 2077 990 2087
rect 121 1890 282 1902
rect 121 1411 136 1890
rect 256 1411 282 1890
rect 916 1467 990 1477
rect 121 1340 282 1411
rect 1161 1340 1183 2323
rect 121 1313 1183 1340
rect 121 1165 233 1313
rect 1058 1280 1183 1313
rect 1291 1280 1315 2323
rect 1991 1922 7491 1932
rect 1991 1731 2084 1922
rect 1991 1721 7491 1731
rect 1412 1572 1574 1580
rect 1406 1570 2248 1572
rect 1406 1496 1412 1570
rect 1574 1562 2248 1570
rect 1574 1502 2196 1562
rect 1574 1496 2248 1502
rect 1406 1492 2248 1496
rect 2454 1562 3538 1572
rect 2506 1502 2970 1562
rect 3022 1502 3486 1562
rect 2454 1492 3538 1502
rect 3744 1562 4828 1572
rect 3796 1502 4260 1562
rect 4312 1502 4776 1562
rect 3744 1492 4828 1502
rect 5034 1562 6118 1572
rect 5086 1502 5550 1562
rect 5602 1502 6066 1562
rect 5034 1492 6118 1502
rect 6324 1562 7408 1572
rect 6376 1502 6840 1562
rect 6892 1502 7356 1562
rect 6324 1492 7408 1502
rect 1412 1486 1574 1492
rect 2712 1446 3280 1456
rect 2764 1386 3228 1446
rect 2712 1376 3280 1386
rect 4002 1446 4570 1456
rect 4054 1386 4518 1446
rect 4002 1376 4570 1386
rect 5292 1446 5860 1456
rect 5344 1386 5808 1446
rect 5292 1376 5860 1386
rect 6582 1446 7150 1456
rect 6634 1386 7098 1446
rect 6582 1376 7150 1386
rect 7356 1446 7408 1492
rect 1058 1165 1315 1280
rect 121 1150 1315 1165
rect 270 894 629 904
rect 270 819 629 829
rect 724 894 1083 904
rect 724 819 1083 829
rect 650 774 702 784
rect 390 449 442 468
rect 650 449 702 698
rect 1311 774 1375 784
rect 1827 774 1891 784
rect 1311 624 1375 634
rect 1575 738 1627 748
rect 2970 775 3022 1376
rect 1827 624 1891 634
rect 2512 722 2564 732
rect 1575 451 1627 598
rect 4260 775 4312 1376
rect 2970 652 3022 662
rect 3802 722 3854 732
rect 1017 449 2003 451
rect 24 441 2003 449
rect 24 439 1017 441
rect 23 307 24 383
rect 2512 338 2564 599
rect 5550 775 5602 1376
rect 4260 652 4312 662
rect 5092 722 5144 732
rect 3802 338 3854 599
rect 6840 775 6892 1376
rect 7356 1063 7408 1386
rect 7356 1014 7667 1063
rect 5550 652 5602 662
rect 6382 723 6434 733
rect 5092 338 5144 599
rect 7421 775 7473 1014
rect 7630 1011 7667 1014
rect 6840 643 6892 652
rect 6963 722 7015 732
rect 6382 344 6434 599
rect 7421 642 7473 652
rect 6963 344 7015 599
rect 6167 338 7713 344
rect 23 306 1017 307
rect 23 303 2003 306
rect 2341 334 7713 338
rect 2341 328 6167 334
rect 2341 303 2514 328
rect 23 239 2514 303
rect -22 234 2514 239
rect -33 228 2514 234
rect -33 80 25 228
rect 2004 189 2514 228
rect 2004 183 6167 189
rect 7521 183 7713 334
rect 2004 80 7713 183
rect -33 70 7713 80
rect -22 36 7713 70
<< via2 >>
rect 304 4979 368 5179
rect 1852 4979 1916 5179
rect 3400 4979 3464 5179
rect 4948 4979 5012 5179
rect 6496 4979 6560 5179
rect 566 4403 622 4603
rect 1598 4403 1654 4603
rect 2114 4403 2170 4603
rect 3146 4403 3202 4603
rect 3662 4403 3718 4603
rect 4694 4403 4750 4603
rect 5210 4403 5266 4603
rect 6242 4403 6298 4603
rect 1078 3498 1142 3698
rect 2626 3498 2690 3698
rect 4174 3498 4238 3698
rect 5722 3498 5786 3698
rect 824 2923 880 3123
rect 1340 2922 1396 3122
rect 2372 2922 2428 3122
rect 2888 2922 2944 3122
rect 3920 2922 3976 3122
rect 4436 2922 4492 3122
rect 5468 2922 5524 3122
rect 5984 2922 6040 3122
rect 916 1477 990 2077
rect 1412 1496 1574 1570
rect 270 829 629 894
rect 724 829 1083 894
rect 1311 634 1375 774
rect 1827 634 1891 774
<< metal3 >>
rect 294 5179 378 5184
rect 294 4979 304 5179
rect 368 4979 378 5179
rect 294 4974 378 4979
rect 1842 5179 1926 5184
rect 1842 4979 1852 5179
rect 1916 4979 1926 5179
rect 1842 4974 1926 4979
rect 3390 5179 3474 5184
rect 3390 4979 3400 5179
rect 3464 4979 3474 5179
rect 3390 4974 3474 4979
rect 4938 5179 5022 5184
rect 4938 4979 4948 5179
rect 5012 4979 5022 5179
rect 4938 4974 5022 4979
rect 6486 5179 6570 5184
rect 6486 4979 6496 5179
rect 6560 4979 6570 5179
rect 6486 4974 6570 4979
rect 556 4603 632 4608
rect 556 4474 566 4603
rect 166 4403 566 4474
rect 622 4474 632 4603
rect 1588 4603 1664 4608
rect 1588 4474 1598 4603
rect 622 4403 1598 4474
rect 1654 4474 1664 4603
rect 2104 4603 2180 4608
rect 2104 4474 2114 4603
rect 1654 4403 2114 4474
rect 2170 4474 2180 4603
rect 3136 4603 3212 4608
rect 3136 4474 3146 4603
rect 2170 4403 3146 4474
rect 3202 4474 3212 4603
rect 3652 4603 3728 4608
rect 3652 4474 3662 4603
rect 3202 4403 3662 4474
rect 3718 4474 3728 4603
rect 4684 4603 4760 4608
rect 4684 4474 4694 4603
rect 3718 4403 4694 4474
rect 4750 4474 4760 4603
rect 5200 4603 5276 4608
rect 5200 4474 5210 4603
rect 4750 4403 5210 4474
rect 5266 4474 5276 4603
rect 6232 4603 6308 4608
rect 6232 4474 6242 4603
rect 5266 4403 6242 4474
rect 6298 4403 6308 4603
rect 166 4400 6308 4403
rect 166 2993 240 4400
rect 556 4398 632 4400
rect 1588 4398 1664 4400
rect 2104 4398 2180 4400
rect 3136 4398 3212 4400
rect 3652 4398 3728 4400
rect 4684 4398 4760 4400
rect 5200 4398 5276 4400
rect 6168 4398 6308 4400
rect 1068 3698 1152 3703
rect 1068 3498 1078 3698
rect 1142 3498 1152 3698
rect 1068 3493 1152 3498
rect 2616 3698 2700 3703
rect 2616 3498 2626 3698
rect 2690 3498 2700 3698
rect 2616 3493 2700 3498
rect 4164 3698 4248 3703
rect 4164 3498 4174 3698
rect 4238 3498 4248 3698
rect 4164 3493 4248 3498
rect 5712 3698 5796 3703
rect 5712 3498 5722 3698
rect 5786 3498 5796 3698
rect 5712 3493 5796 3498
rect 814 3123 890 3128
rect 814 2993 824 3123
rect 166 2923 824 2993
rect 880 2993 890 3123
rect 1330 3122 1406 3127
rect 1330 2993 1340 3122
rect 880 2923 1340 2993
rect 166 2922 1340 2923
rect 1396 2993 1406 3122
rect 2362 3122 2438 3127
rect 2362 2993 2372 3122
rect 1396 2922 2372 2993
rect 2428 2993 2438 3122
rect 2878 3122 2954 3127
rect 2878 2993 2888 3122
rect 2428 2922 2888 2993
rect 2944 2993 2954 3122
rect 3910 3122 3986 3127
rect 3910 2993 3920 3122
rect 2944 2922 3920 2993
rect 3976 2993 3986 3122
rect 4426 3122 4502 3127
rect 4426 2993 4436 3122
rect 3976 2922 4436 2993
rect 4492 2993 4502 3122
rect 5458 3122 5534 3127
rect 5458 2993 5468 3122
rect 4492 2922 5468 2993
rect 5524 2993 5534 3122
rect 5974 3122 6050 3127
rect 5974 2993 5984 3122
rect 5524 2922 5984 2993
rect 6040 2922 6050 3122
rect 166 2917 6050 2922
rect 906 2077 1000 2082
rect 906 1477 916 2077
rect 990 1477 1000 2077
rect 1406 1575 1482 2917
rect 1402 1570 1584 1575
rect 1402 1496 1412 1570
rect 1574 1496 1584 1570
rect 1402 1491 1584 1496
rect 906 1472 1000 1477
rect 260 894 639 899
rect 260 829 270 894
rect 629 829 639 894
rect 260 824 639 829
rect 714 894 1093 899
rect 714 829 724 894
rect 1083 829 1093 894
rect 714 824 1093 829
rect 1301 774 1385 779
rect 1301 634 1311 774
rect 1375 634 1385 774
rect 1301 629 1385 634
rect 1817 774 1901 779
rect 1817 634 1827 774
rect 1891 634 1901 774
rect 1817 629 1901 634
<< via3 >>
rect 304 4979 368 5179
rect 1852 4979 1916 5179
rect 3400 4979 3464 5179
rect 4948 4979 5012 5179
rect 6496 4979 6560 5179
rect 1078 3498 1142 3698
rect 2626 3498 2690 3698
rect 4174 3498 4238 3698
rect 5722 3498 5786 3698
rect 916 1477 990 2077
rect 270 829 629 894
rect 724 829 1083 894
rect 1311 634 1375 774
rect 1827 634 1891 774
<< metal4 >>
rect 20 5179 6561 5180
rect 20 5104 304 5179
rect 20 4449 96 5104
rect 303 4979 304 5104
rect 368 5104 1852 5179
rect 368 4979 369 5104
rect 303 4978 369 4979
rect 1851 4979 1852 5104
rect 1916 5104 3400 5179
rect 1916 4979 1917 5104
rect 1851 4978 1917 4979
rect 3399 4979 3400 5104
rect 3464 5104 4948 5179
rect 3464 4979 3465 5104
rect 3399 4978 3465 4979
rect 4947 4979 4948 5104
rect 5012 5104 6496 5179
rect 5012 4979 5013 5104
rect 4947 4978 5013 4979
rect 6495 4979 6496 5104
rect 6560 4979 6561 5179
rect 6495 4978 6561 4979
rect -168 4372 96 4449
rect -168 899 -92 4372
rect 20 3699 96 4372
rect 20 3698 5787 3699
rect 20 3623 1078 3698
rect 1077 3498 1078 3623
rect 1142 3623 2626 3698
rect 1142 3498 1143 3623
rect 1077 3497 1143 3498
rect 2625 3498 2626 3623
rect 2690 3623 4174 3698
rect 2690 3498 2691 3623
rect 2625 3497 2691 3498
rect 4173 3498 4174 3623
rect 4238 3623 5722 3698
rect 4238 3498 4239 3623
rect 4173 3497 4239 3498
rect 5721 3498 5722 3623
rect 5786 3498 5787 3698
rect 5721 3497 5787 3498
rect 915 2077 991 2078
rect 915 1477 916 2077
rect 990 1548 991 2077
rect 990 1477 1637 1548
rect 915 1472 1637 1477
rect 1571 1080 1637 1472
rect 1310 1004 1892 1080
rect -168 894 1121 899
rect -168 829 270 894
rect 629 829 724 894
rect 1083 829 1121 894
rect -168 826 1121 829
rect 1310 774 1376 1004
rect 1310 634 1311 774
rect 1375 634 1376 774
rect 1310 633 1376 634
rect 1826 774 1892 1004
rect 1826 634 1827 774
rect 1891 634 1892 774
rect 1826 633 1892 634
<< labels >>
rlabel metal2 7711 193 7711 193 7 vcc
port 1 w
rlabel metal2 -51 5514 -51 5514 3 vss
port 2 e
rlabel metal2 7666 1038 7666 1038 7 vref
port 3 w
rlabel metal2 -32 153 -32 153 7 BGR_BJT_stage1_0.vcc
rlabel metal2 -4 5517 -4 5517 7 BGR_BJT_stage1_0.vss
rlabel metal3 1439 2213 1439 2213 5 BGR_BJT_stage1_0.vref0
rlabel metal1 2032 851 2032 851 3 BGR_BJT_stage1_0.vr
flabel locali 607 1733 855 1837 0 FreeSans 400 0 0 0 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter
flabel locali 666 2359 767 2408 0 FreeSans 400 0 0 0 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Collector
flabel locali 643 2209 761 2249 0 FreeSans 400 0 0 0 BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Base
rlabel metal2 2466 257 2466 257 3 BGR_BJT_stage2_0.vcc
rlabel metal2 1992 1848 1992 1848 3 BGR_BJT_stage2_0.vss
rlabel metal2 1961 1528 1961 1528 3 BGR_BJT_stage2_0.vref0
rlabel metal1 2394 848 2394 848 3 BGR_BJT_stage2_0.vr
rlabel metal2 7633 1038 7633 1038 7 BGR_BJT_stage2_0.vref
<< end >>
