magic
tech sky130A
magscale 1 2
timestamp 1741058913
<< pwell >>
rect -201 -702 201 702
<< psubdiff >>
rect -165 632 -69 666
rect 69 632 165 666
rect -165 570 -131 632
rect 131 570 165 632
rect -165 -632 -131 -570
rect 131 -632 165 -570
rect -165 -666 -69 -632
rect 69 -666 165 -632
<< psubdiffcont >>
rect -69 632 69 666
rect -165 -570 -131 570
rect 131 -570 165 570
rect -69 -666 69 -632
<< xpolycontact >>
rect -35 104 35 536
rect -35 -536 35 -104
<< xpolyres >>
rect -35 -104 35 104
<< locali >>
rect -165 632 -69 666
rect 69 632 165 666
rect -165 570 -131 632
rect 131 570 165 632
rect -165 -632 -131 -570
rect 131 -632 165 -570
rect -165 -666 -69 -632
rect 69 -666 165 -632
<< viali >>
rect -19 121 19 518
rect -19 -518 19 -121
<< metal1 >>
rect -25 518 25 530
rect -25 121 -19 518
rect 19 121 25 518
rect -25 109 25 121
rect -25 -121 25 -109
rect -25 -518 -19 -121
rect 19 -518 25 -121
rect -25 -530 25 -518
<< properties >>
string FIXED_BBOX -148 -649 148 649
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.2 m 1 nx 1 wmin 0.350 lmin 0.50 class resistor rho 2000 val 7.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 mult 1
<< end >>
