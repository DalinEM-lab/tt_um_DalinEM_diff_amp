magic
tech sky130A
magscale 1 2
timestamp 1738282926
<< nwell >>
rect -296 -339 296 339
<< pmoslvt >>
rect -100 -120 100 120
<< pdiff >>
rect -158 108 -100 120
rect -158 -108 -146 108
rect -112 -108 -100 108
rect -158 -120 -100 -108
rect 100 108 158 120
rect 100 -108 112 108
rect 146 -108 158 108
rect 100 -120 158 -108
<< pdiffc >>
rect -146 -108 -112 108
rect 112 -108 146 108
<< nsubdiff >>
rect -260 269 -164 303
rect 164 269 260 303
rect -260 207 -226 269
rect 226 207 260 269
rect -260 -269 -226 -207
rect 226 -269 260 -207
rect -260 -303 -164 -269
rect 164 -303 260 -269
<< nsubdiffcont >>
rect -164 269 164 303
rect -260 -207 -226 207
rect 226 -207 260 207
rect -164 -303 164 -269
<< poly >>
rect -100 201 100 217
rect -100 167 -84 201
rect 84 167 100 201
rect -100 120 100 167
rect -100 -167 100 -120
rect -100 -201 -84 -167
rect 84 -201 100 -167
rect -100 -217 100 -201
<< polycont >>
rect -84 167 84 201
rect -84 -201 84 -167
<< locali >>
rect -260 269 -164 303
rect 164 269 260 303
rect -260 207 -226 269
rect 226 207 260 269
rect -100 167 -84 201
rect 84 167 100 201
rect -146 108 -112 124
rect -146 -124 -112 -108
rect 112 108 146 124
rect 112 -124 146 -108
rect -100 -201 -84 -167
rect 84 -201 100 -167
rect -260 -269 -226 -207
rect 226 -269 260 -207
rect -260 -303 -164 -269
rect 164 -303 260 -269
<< viali >>
rect -84 167 84 201
rect -146 -108 -112 108
rect 112 -108 146 108
rect -84 -201 84 -167
<< metal1 >>
rect -96 201 96 207
rect -96 167 -84 201
rect 84 167 96 201
rect -96 161 96 167
rect -152 108 -106 120
rect -152 -108 -146 108
rect -112 -108 -106 108
rect -152 -120 -106 -108
rect 106 108 152 120
rect 106 -108 112 108
rect 146 -108 152 108
rect 106 -120 152 -108
rect -96 -167 96 -161
rect -96 -201 -84 -167
rect 84 -201 96 -167
rect -96 -207 96 -201
<< properties >>
string FIXED_BBOX -243 -286 243 286
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.2 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>
