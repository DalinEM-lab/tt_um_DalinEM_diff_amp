* NGSPICE file created from OTA_stage2_flat.ext - technology: sky130A

.subckt OTA_stage2_flat vcc vss vo vd1 vd2 vb1
X0 a_6817_n2960.t11 vd2.t0 a_7255_n2960.t5 vcc.t3 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X1 a_7255_n2960.t7 vd2.t1 a_6817_n2960.t10 vcc.t2 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X2 vcc.t1 vb1.t0 a_7255_n2960.t0 vcc.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=81200,2916 d=40600,1458
X3 a_14590_n1959.t1 vd1.t0 sky130_fd_pr__cap_mim_m3_1 l=20 w=20
X4 a_7255_n2960.t4 vd1.t1 vo.t4 vcc.t5 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X5 vo.t5 a_6817_n2960.t12 vss.t12 vss.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X6 vo.t3 vd1.t2 a_7255_n2960.t3 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X7 vss.t11 a_6817_n2960.t4 a_6817_n2960.t5 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X8 vo.t2 vd1.t3 a_7255_n2960.t2 vcc.t3 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X9 vss.t10 a_6817_n2960.t13 vo.t6 vss.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X10 a_6817_n2960.t7 a_6817_n2960.t6 vss.t9 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X11 a_14590_n1959.t0 vo.t0 vss.t0 sky130_fd_pr__res_xhigh_po_0p35 l=1
X12 vcc.t9 vb1.t1 a_7255_n2960.t10 vcc.t8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X13 a_7255_n2960.t9 vb1.t2 vcc.t7 vcc.t6 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=81200,2916
X14 a_7255_n2960.t1 vd1.t4 vo.t1 vcc.t2 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X15 a_6817_n2960.t9 vd2.t2 a_7255_n2960.t8 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X16 a_6817_n2960.t3 a_6817_n2960.t2 vss.t8 vss.t7 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X17 a_7255_n2960.t11 vb1.t3 vcc.t11 vcc.t10 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X18 a_7255_n2960.t6 vd2.t3 a_6817_n2960.t8 vcc.t5 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X19 vss.t6 a_6817_n2960.t14 vo.t7 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X20 vss.t4 a_6817_n2960.t0 a_6817_n2960.t1 vss.t3 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X21 vo.t8 a_6817_n2960.t15 vss.t2 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
R0 vd2.n0 vd2.t0 122.688
R1 vd2.n1 vd2.t2 122.213
R2 vd2.n0 vd2.t1 122.213
R3 vd2.n2 vd2.t3 121.831
R4 vd2 vd2.n2 1.1155
R5 vd2.n1 vd2.n0 0.548
R6 vd2.n2 vd2.n1 0.238
R7 a_7255_n2960.n0 a_7255_n2960.t9 36.4777
R8 a_7255_n2960.n0 a_7255_n2960.t0 35.4327
R9 a_7255_n2960.n0 a_7255_n2960.n4 31.3519
R10 a_7255_n2960.n7 a_7255_n2960.n6 18.3035
R11 a_7255_n2960.n3 a_7255_n2960.n2 18.303
R12 a_7255_n2960.n8 a_7255_n2960.n7 17.2098
R13 a_7255_n2960.n3 a_7255_n2960.n1 17.208
R14 a_7255_n2960.n5 a_7255_n2960.n3 8.938
R15 a_7255_n2960.n4 a_7255_n2960.t10 4.08121
R16 a_7255_n2960.n4 a_7255_n2960.t11 4.08121
R17 a_7255_n2960.n5 a_7255_n2960.n0 3.2905
R18 a_7255_n2960.n7 a_7255_n2960.n5 3.05142
R19 a_7255_n2960.n2 a_7255_n2960.t8 1.90483
R20 a_7255_n2960.n2 a_7255_n2960.t4 1.90483
R21 a_7255_n2960.n1 a_7255_n2960.t2 1.90483
R22 a_7255_n2960.n1 a_7255_n2960.t7 1.90483
R23 a_7255_n2960.n6 a_7255_n2960.t3 1.90483
R24 a_7255_n2960.n6 a_7255_n2960.t6 1.90483
R25 a_7255_n2960.n8 a_7255_n2960.t5 1.90483
R26 a_7255_n2960.t1 a_7255_n2960.n8 1.90483
R27 a_6817_n2960.n3 a_6817_n2960.t3 60.3532
R28 a_6817_n2960.n10 a_6817_n2960.t1 60.3532
R29 a_6817_n2960.n15 a_6817_n2960.n14 48.5755
R30 a_6817_n2960.n0 a_6817_n2960.t8 19.1315
R31 a_6817_n2960.t11 a_6817_n2960.n0 18.308
R32 a_6817_n2960.n0 a_6817_n2960.n1 16.2734
R33 a_6817_n2960.n12 a_6817_n2960.n11 14.6534
R34 a_6817_n2960.n14 a_6817_n2960.t5 11.6005
R35 a_6817_n2960.n14 a_6817_n2960.t7 11.6005
R36 a_6817_n2960.n10 a_6817_n2960.n2 11.2227
R37 a_6817_n2960.n16 a_6817_n2960.n15 8.08817
R38 a_6817_n2960.n3 a_6817_n2960.n2 7.9105
R39 a_6817_n2960.n4 a_6817_n2960.t2 3.58326
R40 a_6817_n2960.n6 a_6817_n2960.t14 3.58326
R41 a_6817_n2960.n8 a_6817_n2960.t15 3.58326
R42 a_6817_n2960.n9 a_6817_n2960.t0 3.58326
R43 a_6817_n2960.n4 a_6817_n2960.t12 3.58267
R44 a_6817_n2960.n6 a_6817_n2960.t4 3.58267
R45 a_6817_n2960.n8 a_6817_n2960.t6 3.58267
R46 a_6817_n2960.n9 a_6817_n2960.t13 3.58267
R47 a_6817_n2960.n13 a_6817_n2960.n12 3.54985
R48 a_6817_n2960.n0 a_6817_n2960.n16 2.67636
R49 a_6817_n2960.n16 a_6817_n2960.n2 2.10354
R50 a_6817_n2960.n1 a_6817_n2960.t10 1.90483
R51 a_6817_n2960.n1 a_6817_n2960.t9 1.90483
R52 a_6817_n2960.n7 a_6817_n2960.n5 1.69798
R53 a_6817_n2960.n11 a_6817_n2960.n9 1.61224
R54 a_6817_n2960.n12 a_6817_n2960.n8 1.61224
R55 a_6817_n2960.n7 a_6817_n2960.n6 1.61224
R56 a_6817_n2960.n5 a_6817_n2960.n4 1.61224
R57 a_6817_n2960.n11 a_6817_n2960.n10 0.995611
R58 a_6817_n2960.n5 a_6817_n2960.n3 0.96988
R59 a_6817_n2960.n15 a_6817_n2960.n13 0.793374
R60 a_6817_n2960.n13 a_6817_n2960.n7 0.432312
R61 vcc.n45 vcc.n2 17565.9
R62 vcc.n45 vcc.n3 17565.9
R63 vcc.n43 vcc.n3 17562.4
R64 vcc.n43 vcc.n2 17562.4
R65 vcc.n29 vcc.n13 6349.41
R66 vcc.n29 vcc.n14 6349.41
R67 vcc.n27 vcc.n13 6349.41
R68 vcc.n27 vcc.n14 6349.41
R69 vcc.t8 vcc.t6 216.05
R70 vcc.t10 vcc.t0 216.05
R71 vcc.n47 vcc.n1 209.422
R72 vcc.t6 vcc.n13 174.992
R73 vcc.t0 vcc.n14 174.992
R74 vcc.n46 vcc.n0 157.375
R75 vcc.n37 vcc.n36 116.722
R76 vcc.n6 vcc.n5 115.912
R77 vcc.n5 vcc.n0 108.909
R78 vcc.n28 vcc.t8 108.025
R79 vcc.n28 vcc.t10 108.025
R80 vcc.n42 vcc.n41 87.9664
R81 vcc.n41 vcc.n6 87.7954
R82 vcc.n17 vcc.n16 71.8902
R83 vcc.t3 vcc.n2 71.3347
R84 vcc.n26 vcc.n15 70.7824
R85 vcc.n33 vcc.n8 65.6211
R86 vcc.t5 vcc.n3 60.8049
R87 vcc.n9 vcc.n1 55.3321
R88 vcc.t2 vcc.t3 53.6285
R89 vcc.t4 vcc.t5 53.6285
R90 vcc.n30 vcc.n12 50.9389
R91 vcc.n20 vcc.n18 32.1789
R92 vcc.n44 vcc.t4 32.0794
R93 vcc.n20 vcc.n19 32.0774
R94 vcc.n36 vcc.n8 30.7043
R95 vcc.n31 vcc.n30 30.0503
R96 vcc.n31 vcc.n11 29.6052
R97 vcc.n44 vcc.t2 21.5497
R98 vcc.n38 vcc.n37 9.34567
R99 vcc.n25 vcc.n24 9.3005
R100 vcc.n34 vcc.n33 9.3005
R101 vcc.n41 vcc.n40 9.3005
R102 vcc.n16 vcc.n14 8.04398
R103 vcc.n15 vcc.n13 8.04398
R104 vcc.n27 vcc.n26 7.11588
R105 vcc.n28 vcc.n27 7.11588
R106 vcc.n30 vcc.n29 7.11588
R107 vcc.n29 vcc.n28 7.11588
R108 vcc.n9 vcc.n8 6.56253
R109 vcc.n43 vcc.n42 5.44168
R110 vcc.n44 vcc.n43 5.44168
R111 vcc.n46 vcc.n45 5.44168
R112 vcc.n45 vcc.n44 5.44168
R113 vcc.n26 vcc.n25 4.82369
R114 vcc.n15 vcc.n12 4.48345
R115 vcc.n37 vcc.n4 4.42232
R116 vcc.n18 vcc.t7 4.08121
R117 vcc.n18 vcc.t9 4.08121
R118 vcc.n19 vcc.t11 4.08121
R119 vcc.n19 vcc.t1 4.08121
R120 vcc.n25 vcc.n17 1.94833
R121 vcc.n38 vcc.n7 1.87667
R122 vcc.n42 vcc.n4 1.86232
R123 vcc.n2 vcc.n1 1.66717
R124 vcc.n5 vcc.n3 1.66717
R125 vcc.n32 vcc.n31 1.6211
R126 vcc.n47 vcc.n46 1.20392
R127 vcc.n16 vcc.n11 1.19816
R128 vcc.n35 vcc.n34 0.985286
R129 vcc.n40 vcc.n39 0.96321
R130 vcc.n23 vcc.n22 0.928261
R131 vcc.n36 vcc.n35 0.875256
R132 vcc.n21 vcc.n12 0.872492
R133 vcc.n35 vcc.n9 0.862026
R134 vcc.n40 vcc.n7 0.758322
R135 vcc.n48 vcc.n0 0.730191
R136 vcc.n22 vcc.n21 0.445398
R137 vcc.n48 vcc.n47 0.428528
R138 vcc.n7 vcc.n6 0.342518
R139 vcc vcc.n48 0.339989
R140 vcc.n33 vcc.n32 0.137839
R141 vcc.n22 vcc.n11 0.129667
R142 vcc.n39 vcc.n4 0.129667
R143 vcc.n23 vcc.n17 0.103833
R144 vcc.n24 vcc.n20 0.047375
R145 vcc.n32 vcc.n10 0.0341957
R146 vcc.n24 vcc.n23 0.0216694
R147 vcc.n21 vcc.n10 0.020648
R148 vcc.n34 vcc.n10 0.00255592
R149 vcc.n39 vcc.n38 0.00155302
R150 vb1.n0 vb1.t0 68.1062
R151 vb1.n0 vb1.t3 67.5138
R152 vb1.n1 vb1.t1 67.5138
R153 vb1.n2 vb1.t2 67.5138
R154 vb1 vb1.n2 8.86177
R155 vb1.n1 vb1.n0 0.603761
R156 vb1.n2 vb1.n1 0.557565
R157 a_14590_n1959.t0 a_14590_n1959.t1 53.247
R158 vd1.n2 vd1.t2 122.216
R159 vd1.n1 vd1.t4 122.216
R160 vd1.n3 vd1.t1 121.828
R161 vd1.n0 vd1.t3 121.828
R162 vd1.n0 vd1.t0 5.15117
R163 vd1.n3 vd1.n2 0.858
R164 vd1 vd1.n3 0.8055
R165 vd1.n2 vd1.n1 0.548
R166 vd1.n1 vd1.n0 0.238
R167 vo.n3 vo.t6 72.7606
R168 vo.n4 vo.t5 71.6732
R169 vo vo.n6 62.2269
R170 vo.n5 vo.t0 52.9855
R171 vo.n0 vo.t4 19.4751
R172 vo.n0 vo.t2 18.6511
R173 vo.n2 vo.n1 15.6099
R174 vo.n6 vo.t7 11.6005
R175 vo.n6 vo.t8 11.6005
R176 vo.n4 vo.n3 2.48505
R177 vo.n1 vo.t1 1.90483
R178 vo.n1 vo.t3 1.90483
R179 vo.n2 vo.n0 1.32214
R180 vo.n3 vo.n2 1.28407
R181 vo vo.n5 0.361755
R182 vo.n5 vo.n4 0.00787255
R183 vss.n45 vss.n44 874968
R184 vss.n21 vss.n10 27614.8
R185 vss.n46 vss.n10 27609
R186 vss.n21 vss.n11 27609
R187 vss.n46 vss.n11 27603.2
R188 vss.n19 vss.n13 4403.53
R189 vss.n19 vss.n14 4403.53
R190 vss.n42 vss.n13 4403.53
R191 vss.n42 vss.n14 4403.53
R192 vss.t7 vss.t5 4074.72
R193 vss.t1 vss.t3 3478.61
R194 vss.n45 vss.t3 2794.88
R195 vss.t5 vss.n12 1000.75
R196 vss.n43 vss.t7 959.708
R197 vss.n48 vss.n8 903.91
R198 vss.n44 vss.t1 610.412
R199 vss.n44 vss.n12 532.535
R200 vss.n16 vss.n14 292.5
R201 vss.n14 vss.t0 292.5
R202 vss.n15 vss.n13 292.5
R203 vss.n13 vss.t0 292.5
R204 vss.n36 vss.n35 262.366
R205 vss.n26 vss.n24 252.304
R206 vss.n22 vss.n17 223.468
R207 vss.n20 vss.t0 169.495
R208 vss.n50 vss.n7 169.446
R209 vss.n21 vss.n20 165.347
R210 vss.n44 vss.n43 106.507
R211 vss.n18 vss.n15 68.9197
R212 vss.n23 vss.n22 68.8547
R213 vss.n18 vss.n16 67.4522
R214 vss.n41 vss.n15 67.2825
R215 vss.n44 vss.t0 62.9885
R216 vss.n30 vss.n29 56.2007
R217 vss.n5 vss.n4 55.1712
R218 vss.n31 vss.n28 54.0035
R219 vss.n2 vss.n1 53.9338
R220 vss.n41 vss.n40 51.5266
R221 vss.n47 vss.n9 39.7638
R222 vss.n50 vss.n49 39.511
R223 vss.n39 vss.n23 37.2591
R224 vss.n40 vss.n39 36.6884
R225 vss.n19 vss.n18 36.563
R226 vss.n20 vss.n19 36.563
R227 vss.n42 vss.n41 36.563
R228 vss.n43 vss.n42 36.563
R229 vss.n22 vss.n21 32.5005
R230 vss.n47 vss.n46 32.5005
R231 vss.n46 vss.n45 32.5005
R232 vss.n36 vss.n26 15.5385
R233 vss.n40 vss.n16 14.2889
R234 vss.n4 vss.t8 11.6005
R235 vss.n4 vss.t6 11.6005
R236 vss.n1 vss.t2 11.6005
R237 vss.n1 vss.t4 11.6005
R238 vss.n28 vss.t9 11.6005
R239 vss.n28 vss.t10 11.6005
R240 vss.n29 vss.t12 11.6005
R241 vss.n29 vss.t11 11.6005
R242 vss.n17 vss.n7 10.5495
R243 vss.n38 vss.n24 9.35616
R244 vss.n33 vss.n8 9.30287
R245 vss.n51 vss.n50 9.3005
R246 vss.n35 vss.n34 9.3005
R247 vss.n17 vss.n11 4.8755
R248 vss.n12 vss.n11 4.8755
R249 vss.n26 vss.n10 4.8755
R250 vss.n12 vss.n10 4.8755
R251 vss.n52 vss.n51 4.5005
R252 vss.n38 vss.n37 4.1842
R253 vss.n27 vss.n25 4.11666
R254 vss.n35 vss.n9 3.76521
R255 vss.n51 vss.n6 2.34664
R256 vss.n33 vss.n32 2.29449
R257 vss.n32 vss.n31 2.11733
R258 vss.n31 vss.n30 1.74237
R259 vss.n49 vss.n48 1.30961
R260 vss.n52 vss.n2 1.21619
R261 vss.n48 vss.n47 1.06085
R262 vss.n5 vss.n2 0.995892
R263 vss.n39 vss.n38 0.874635
R264 vss.n9 vss.n8 0.684992
R265 vss.n32 vss.n0 0.55067
R266 vss.n53 vss.n0 0.497949
R267 vss.n27 vss.n3 0.484781
R268 vss.n51 vss.n3 0.446546
R269 vss.n49 vss.n3 0.32741
R270 vss.n24 vss.n23 0.205848
R271 vss.n3 vss.n0 0.1255
R272 vss.n37 vss.n36 0.0850455
R273 vss vss.n53 0.0796284
R274 vss.n34 vss.n27 0.0386737
R275 vss.n30 vss.n25 0.0370854
R276 vss.n37 vss.n25 0.0287609
R277 vss.n7 vss.n6 0.0286818
R278 vss.n53 vss.n52 0.0274495
R279 vss.n6 vss.n5 0.0126951
R280 vss.n34 vss.n33 0.0028696
C0 vo vb1 0.211041f
C1 vo vd2 0.970649f
C2 vo vd1 6.13476f
C3 vd1 vd2 2.47175f
C4 vcc vb1 7.65782f
C5 vo vcc 3.91529f
C6 vcc vd2 3.74243f
C7 vcc vd1 4.15541f
C8 vb1 vss 3.782027f
C9 vo vss 12.790721f
C10 vd2 vss 2.220361f
C11 vd1 vss 13.139122f
C12 vcc vss 92.16464f
C13 vo.t0 vss 0.10054f
C14 vo.t2 vss 0.737802f
C15 vo.t4 vss 0.820006f
C16 vo.n0 vss 4.30737f
C17 vo.t1 vss 0.155122f
C18 vo.t3 vss 0.155122f
C19 vo.n1 vss 0.430854f
C20 vo.n2 vss 2.50131f
C21 vo.t6 vss 0.084338f
C22 vo.n3 vss 2.47769f
C23 vo.t5 vss 0.076084f
C24 vo.n4 vss 1.14326f
C25 vo.n5 vss 0.791679f
C26 vo.t7 vss 0.015512f
C27 vo.t8 vss 0.015512f
C28 vo.n6 vss 0.091281f
C29 vd1.t0 vss 37.0822f
C30 vd1.t3 vss 1.57149f
C31 vd1.n0 vss 2.9213f
C32 vd1.t4 vss 1.5819f
C33 vd1.n1 vss 2.61695f
C34 vd1.t2 vss 1.5819f
C35 vd1.n2 vss 2.6691f
C36 vd1.t1 vss 1.57149f
C37 vd1.n3 vss 2.63577f
C38 a_14590_n1959.t1 vss 35.8635f
C39 a_14590_n1959.t0 vss 0.036479f
C40 vb1.t0 vss 0.989256f
C41 vb1.t3 vss 0.97562f
C42 vb1.n0 vss 3.14441f
C43 vb1.t1 vss 0.97562f
C44 vb1.n1 vss 1.5897f
C45 vb1.t2 vss 0.97562f
C46 vb1.n2 vss 1.89715f
C47 vcc.n0 vss 0.989659f
C48 vcc.n1 vss 0.528892f
C49 vcc.n2 vss 2.30815f
C50 vcc.n3 vss 1.93657f
C51 vcc.t3 vss 2.73333f
C52 vcc.t2 vss 1.63463f
C53 vcc.n4 vss 0.004585f
C54 vcc.n5 vss 0.329991f
C55 vcc.n6 vss 0.651465f
C56 vcc.n7 vss 0.25087f
C57 vcc.n8 vss 0.532263f
C58 vcc.n9 vss 0.174929f
C59 vcc.n10 vss 0.005633f
C60 vcc.n11 vss 0.096576f
C61 vcc.n12 vss 1.34225f
C62 vcc.n13 vss 0.300507f
C63 vcc.n14 vss 0.300507f
C64 vcc.t6 vss 0.479749f
C65 vcc.t8 vss 0.395419f
C66 vcc.n15 vss 0.327455f
C67 vcc.n16 vss 0.22564f
C68 vcc.n17 vss 0.186481f
C69 vcc.t7 vss 0.013931f
C70 vcc.t9 vss 0.013931f
C71 vcc.n18 vss 0.036186f
C72 vcc.t11 vss 0.013931f
C73 vcc.t1 vss 0.013931f
C74 vcc.n19 vss 0.035519f
C75 vcc.n20 vss 0.568352f
C76 vcc.n21 vss 0.965513f
C77 vcc.n22 vss 0.237643f
C78 vcc.n23 vss 0.168971f
C79 vcc.n24 vss 0.181249f
C80 vcc.n25 vss 0.013826f
C81 vcc.n26 vss 0.204426f
C82 vcc.n27 vss 0.042349f
C83 vcc.t0 vss 0.479749f
C84 vcc.t10 vss 0.395419f
C85 vcc.n28 vss 0.263613f
C86 vcc.n29 vss 0.042349f
C87 vcc.n30 vss 0.492466f
C88 vcc.n31 vss 0.277178f
C89 vcc.n32 vss 0.010233f
C90 vcc.n33 vss 0.382785f
C91 vcc.n34 vss 0.250339f
C92 vcc.n35 vss 0.384102f
C93 vcc.n36 vss 0.420245f
C94 vcc.n37 vss 0.126285f
C95 vcc.n38 vss 0.417024f
C96 vcc.n39 vss 0.067985f
C97 vcc.n40 vss 0.166501f
C98 vcc.n41 vss 0.212215f
C99 vcc.n42 vss 0.066433f
C100 vcc.n43 vss 0.116705f
C101 vcc.t5 vss 2.50324f
C102 vcc.t4 vss 1.86358f
C103 vcc.n44 vss 1.16607f
C104 vcc.n45 vss 0.116728f
C105 vcc.n46 vss 0.24377f
C106 vcc.n47 vss 0.918709f
C107 vcc.n48 vss 0.294637f
C108 a_6817_n2960.n0 vss 1.84569f
C109 a_6817_n2960.t10 vss 0.04377f
C110 a_6817_n2960.t9 vss 0.04377f
C111 a_6817_n2960.n1 vss 0.13799f
C112 a_6817_n2960.n2 vss 1.02544f
C113 a_6817_n2960.t3 vss 0.015448f
C114 a_6817_n2960.n3 vss 0.072402f
C115 a_6817_n2960.t2 vss 0.608715f
C116 a_6817_n2960.t12 vss 0.608712f
C117 a_6817_n2960.n4 vss 0.226883f
C118 a_6817_n2960.n5 vss 1.60678f
C119 a_6817_n2960.t14 vss 0.608715f
C120 a_6817_n2960.t4 vss 0.608712f
C121 a_6817_n2960.n6 vss 0.226883f
C122 a_6817_n2960.n7 vss 1.58469f
C123 a_6817_n2960.t15 vss 0.608715f
C124 a_6817_n2960.t6 vss 0.608712f
C125 a_6817_n2960.n8 vss 0.226883f
C126 a_6817_n2960.t0 vss 0.608715f
C127 a_6817_n2960.t13 vss 0.608712f
C128 a_6817_n2960.n9 vss 0.226883f
C129 a_6817_n2960.t1 vss 0.015448f
C130 a_6817_n2960.n10 vss 0.20036f
C131 a_6817_n2960.n11 vss 1.61012f
C132 a_6817_n2960.n12 vss 1.62999f
C133 a_6817_n2960.n13 vss 0.103003f
C134 a_6817_n2960.t5 vss 0.004377f
C135 a_6817_n2960.t7 vss 0.004377f
C136 a_6817_n2960.n14 vss 0.009258f
C137 a_6817_n2960.n15 vss 0.033706f
C138 a_6817_n2960.n16 vss 0.615675f
C139 a_6817_n2960.t8 vss 0.22076f
C140 a_6817_n2960.t11 vss 0.199702f
C141 a_7255_n2960.n0 vss 3.46131f
C142 a_7255_n2960.t5 vss 0.215884f
C143 a_7255_n2960.t2 vss 0.215884f
C144 a_7255_n2960.t7 vss 0.215884f
C145 a_7255_n2960.n1 vss 0.668091f
C146 a_7255_n2960.t8 vss 0.215884f
C147 a_7255_n2960.t4 vss 0.215884f
C148 a_7255_n2960.n2 vss 0.75835f
C149 a_7255_n2960.n3 vss 4.70225f
C150 a_7255_n2960.t0 vss 0.39757f
C151 a_7255_n2960.t10 vss 0.100746f
C152 a_7255_n2960.t11 vss 0.100746f
C153 a_7255_n2960.n4 vss 0.234713f
C154 a_7255_n2960.t9 vss 0.425266f
C155 a_7255_n2960.n5 vss 2.87401f
C156 a_7255_n2960.t3 vss 0.215884f
C157 a_7255_n2960.t6 vss 0.215884f
C158 a_7255_n2960.n6 vss 0.758372f
C159 a_7255_n2960.n7 vss 3.52329f
C160 a_7255_n2960.n8 vss 0.668219f
C161 a_7255_n2960.t1 vss 0.215884f
C162 vd2.t0 vss 1.68308f
C163 vd2.t1 vss 1.67463f
C164 vd2.n0 vss 5.57114f
C165 vd2.t2 vss 1.67463f
C166 vd2.n1 vss 2.77009f
C167 vd2.t3 vss 1.66375f
C168 vd2.n2 vss 2.76316f
.ends

