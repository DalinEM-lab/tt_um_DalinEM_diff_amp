magic
tech sky130A
magscale 1 2
timestamp 1740519234
<< nwell >>
rect 6472 -3262 9085 4497
rect 11508 -3133 13514 -1295
<< pwell >>
rect 14424 -2725 14826 -1361
<< pmos >>
rect 11704 -2914 12064 -1514
rect 12122 -2914 12482 -1514
rect 12540 -2914 12900 -1514
rect 12958 -2914 13318 -1514
<< pmoslvt >>
rect 6875 1017 7255 4017
rect 7313 1017 7693 4017
rect 7751 1017 8131 4017
rect 8189 1017 8569 4017
rect 6875 -2960 7255 40
rect 7313 -2960 7693 40
rect 7751 -2960 8131 40
rect 8189 -2960 8569 40
<< nmoslvt >>
rect 6885 -4286 8765 -3986
rect 8823 -4286 10703 -3986
rect 10761 -4286 12641 -3986
rect 12699 -4286 14579 -3986
rect 6885 -4696 8765 -4396
rect 8823 -4696 10703 -4396
rect 10761 -4696 12641 -4396
rect 12699 -4696 14579 -4396
<< ndiff >>
rect 6827 -3998 6885 -3986
rect 6827 -4274 6839 -3998
rect 6873 -4274 6885 -3998
rect 6827 -4286 6885 -4274
rect 8765 -3998 8823 -3986
rect 8765 -4274 8777 -3998
rect 8811 -4274 8823 -3998
rect 8765 -4286 8823 -4274
rect 10703 -3998 10761 -3986
rect 10703 -4274 10715 -3998
rect 10749 -4274 10761 -3998
rect 10703 -4286 10761 -4274
rect 12641 -3998 12699 -3986
rect 12641 -4274 12653 -3998
rect 12687 -4274 12699 -3998
rect 12641 -4286 12699 -4274
rect 14579 -3998 14637 -3986
rect 14579 -4274 14591 -3998
rect 14625 -4274 14637 -3998
rect 14579 -4286 14637 -4274
rect 6827 -4408 6885 -4396
rect 6827 -4684 6839 -4408
rect 6873 -4684 6885 -4408
rect 6827 -4696 6885 -4684
rect 8765 -4408 8823 -4396
rect 8765 -4684 8777 -4408
rect 8811 -4684 8823 -4408
rect 8765 -4696 8823 -4684
rect 10703 -4408 10761 -4396
rect 10703 -4684 10715 -4408
rect 10749 -4684 10761 -4408
rect 10703 -4696 10761 -4684
rect 12641 -4408 12699 -4396
rect 12641 -4684 12653 -4408
rect 12687 -4684 12699 -4408
rect 12641 -4696 12699 -4684
rect 14579 -4408 14637 -4396
rect 14579 -4684 14591 -4408
rect 14625 -4684 14637 -4408
rect 14579 -4696 14637 -4684
<< pdiff >>
rect 6817 4005 6875 4017
rect 6817 1029 6829 4005
rect 6863 1029 6875 4005
rect 6817 1017 6875 1029
rect 7255 4005 7313 4017
rect 7255 1029 7267 4005
rect 7301 1029 7313 4005
rect 7255 1017 7313 1029
rect 7693 4005 7751 4017
rect 7693 1029 7705 4005
rect 7739 1029 7751 4005
rect 7693 1017 7751 1029
rect 8131 4005 8189 4017
rect 8131 1029 8143 4005
rect 8177 1029 8189 4005
rect 8131 1017 8189 1029
rect 8569 4005 8627 4017
rect 8569 1029 8581 4005
rect 8615 1029 8627 4005
rect 8569 1017 8627 1029
rect 6817 28 6875 40
rect 6817 -2948 6829 28
rect 6863 -2948 6875 28
rect 6817 -2960 6875 -2948
rect 7255 28 7313 40
rect 7255 -2948 7267 28
rect 7301 -2948 7313 28
rect 7255 -2960 7313 -2948
rect 7693 28 7751 40
rect 7693 -2948 7705 28
rect 7739 -2948 7751 28
rect 7693 -2960 7751 -2948
rect 8131 28 8189 40
rect 8131 -2948 8143 28
rect 8177 -2948 8189 28
rect 8131 -2960 8189 -2948
rect 8569 28 8627 40
rect 8569 -2948 8581 28
rect 8615 -2948 8627 28
rect 8569 -2960 8627 -2948
rect 11646 -1526 11704 -1514
rect 11646 -2902 11658 -1526
rect 11692 -2902 11704 -1526
rect 11646 -2914 11704 -2902
rect 12064 -1526 12122 -1514
rect 12064 -2902 12076 -1526
rect 12110 -2902 12122 -1526
rect 12064 -2914 12122 -2902
rect 12482 -1526 12540 -1514
rect 12482 -2902 12494 -1526
rect 12528 -2902 12540 -1526
rect 12482 -2914 12540 -2902
rect 12900 -1526 12958 -1514
rect 12900 -2902 12912 -1526
rect 12946 -2902 12958 -1526
rect 12900 -2914 12958 -2902
rect 13318 -1526 13376 -1514
rect 13318 -2902 13330 -1526
rect 13364 -2902 13376 -1526
rect 13318 -2914 13376 -2902
<< ndiffc >>
rect 6839 -4274 6873 -3998
rect 8777 -4274 8811 -3998
rect 10715 -4274 10749 -3998
rect 12653 -4274 12687 -3998
rect 14591 -4274 14625 -3998
rect 6839 -4684 6873 -4408
rect 8777 -4684 8811 -4408
rect 10715 -4684 10749 -4408
rect 12653 -4684 12687 -4408
rect 14591 -4684 14625 -4408
<< pdiffc >>
rect 6829 1029 6863 4005
rect 7267 1029 7301 4005
rect 7705 1029 7739 4005
rect 8143 1029 8177 4005
rect 8581 1029 8615 4005
rect 6829 -2948 6863 28
rect 7267 -2948 7301 28
rect 7705 -2948 7739 28
rect 8143 -2948 8177 28
rect 8581 -2948 8615 28
rect 11658 -2902 11692 -1526
rect 12076 -2902 12110 -1526
rect 12494 -2902 12528 -1526
rect 12912 -2902 12946 -1526
rect 13330 -2902 13364 -1526
<< psubdiff >>
rect 14460 -1431 14556 -1397
rect 14694 -1431 14790 -1397
rect 14460 -1493 14494 -1431
rect 14756 -1493 14790 -1431
rect 14460 -2655 14494 -2593
rect 14756 -2655 14790 -2593
rect 14460 -2689 14556 -2655
rect 14694 -2689 14790 -2655
rect 6617 -3656 6677 -3622
rect 14846 -3656 14906 -3622
rect 6617 -3682 6651 -3656
rect 14872 -3682 14906 -3656
rect 6617 -4931 6651 -4905
rect 14872 -4931 14906 -4905
rect 6617 -4965 6677 -4931
rect 14846 -4965 14906 -4931
<< nsubdiff >>
rect 6565 4397 6625 4431
rect 8905 4397 8965 4431
rect 6565 4371 6599 4397
rect 8931 4371 8965 4397
rect 6565 -3190 6599 -3164
rect 11544 -1365 11640 -1331
rect 13382 -1365 13478 -1331
rect 11544 -1427 11578 -1365
rect 13444 -1427 13478 -1365
rect 11544 -3063 11578 -3001
rect 13444 -3063 13478 -3001
rect 11544 -3097 11640 -3063
rect 13382 -3097 13478 -3063
rect 8931 -3190 8965 -3164
rect 6565 -3224 6625 -3190
rect 8905 -3224 8965 -3190
<< psubdiffcont >>
rect 14556 -1431 14694 -1397
rect 14460 -2593 14494 -1493
rect 14756 -2593 14790 -1493
rect 14556 -2689 14694 -2655
rect 6677 -3656 14846 -3622
rect 6617 -4905 6651 -3682
rect 14872 -4905 14906 -3682
rect 6677 -4965 14846 -4931
<< nsubdiffcont >>
rect 6625 4397 8905 4431
rect 6565 -3164 6599 4371
rect 8931 -3164 8965 4371
rect 11640 -1365 13382 -1331
rect 11544 -3001 11578 -1427
rect 13444 -3001 13478 -1427
rect 11640 -3097 13382 -3063
rect 6625 -3224 8905 -3190
<< poly >>
rect 6875 4098 7255 4114
rect 6875 4064 6891 4098
rect 7239 4064 7255 4098
rect 6875 4017 7255 4064
rect 7313 4098 7693 4114
rect 7313 4064 7329 4098
rect 7677 4064 7693 4098
rect 7313 4017 7693 4064
rect 7751 4098 8131 4114
rect 7751 4064 7767 4098
rect 8115 4064 8131 4098
rect 7751 4017 8131 4064
rect 8189 4098 8569 4114
rect 8189 4064 8205 4098
rect 8553 4064 8569 4098
rect 8189 4017 8569 4064
rect 6875 970 7255 1017
rect 6875 936 6891 970
rect 7239 936 7255 970
rect 6875 920 7255 936
rect 7313 970 7693 1017
rect 7313 936 7329 970
rect 7677 936 7693 970
rect 7313 920 7693 936
rect 7751 970 8131 1017
rect 7751 936 7767 970
rect 8115 936 8131 970
rect 7751 920 8131 936
rect 8189 970 8569 1017
rect 8189 936 8205 970
rect 8553 936 8569 970
rect 8189 920 8569 936
rect 6875 121 7255 137
rect 6875 87 6891 121
rect 7239 87 7255 121
rect 6875 40 7255 87
rect 7313 121 7693 137
rect 7313 87 7329 121
rect 7677 87 7693 121
rect 7313 40 7693 87
rect 7751 121 8131 137
rect 7751 87 7767 121
rect 8115 87 8131 121
rect 7751 40 8131 87
rect 8189 121 8569 137
rect 8189 87 8205 121
rect 8553 87 8569 121
rect 8189 40 8569 87
rect 6875 -3007 7255 -2960
rect 6875 -3041 6891 -3007
rect 7239 -3041 7255 -3007
rect 6875 -3057 7255 -3041
rect 7313 -3007 7693 -2960
rect 7313 -3041 7329 -3007
rect 7677 -3041 7693 -3007
rect 7313 -3057 7693 -3041
rect 7751 -3007 8131 -2960
rect 7751 -3041 7767 -3007
rect 8115 -3041 8131 -3007
rect 7751 -3057 8131 -3041
rect 8189 -3007 8569 -2960
rect 8189 -3041 8205 -3007
rect 8553 -3041 8569 -3007
rect 8189 -3057 8569 -3041
rect 11704 -1433 12064 -1417
rect 11704 -1467 11720 -1433
rect 12048 -1467 12064 -1433
rect 11704 -1514 12064 -1467
rect 12122 -1433 12482 -1417
rect 12122 -1467 12138 -1433
rect 12466 -1467 12482 -1433
rect 12122 -1514 12482 -1467
rect 12540 -1433 12900 -1417
rect 12540 -1467 12556 -1433
rect 12884 -1467 12900 -1433
rect 12540 -1514 12900 -1467
rect 12958 -1433 13318 -1417
rect 12958 -1467 12974 -1433
rect 13302 -1467 13318 -1433
rect 12958 -1514 13318 -1467
rect 11704 -2961 12064 -2914
rect 11704 -2995 11720 -2961
rect 12048 -2995 12064 -2961
rect 11704 -3011 12064 -2995
rect 12122 -2961 12482 -2914
rect 12122 -2995 12138 -2961
rect 12466 -2995 12482 -2961
rect 12122 -3011 12482 -2995
rect 12540 -2961 12900 -2914
rect 12540 -2995 12556 -2961
rect 12884 -2995 12900 -2961
rect 12540 -3011 12900 -2995
rect 12958 -2961 13318 -2914
rect 12958 -2995 12974 -2961
rect 13302 -2995 13318 -2961
rect 12958 -3011 13318 -2995
rect 6885 -3914 8765 -3898
rect 6885 -3948 6901 -3914
rect 8749 -3948 8765 -3914
rect 6885 -3986 8765 -3948
rect 8823 -3914 10703 -3898
rect 8823 -3948 8839 -3914
rect 10687 -3948 10703 -3914
rect 8823 -3986 10703 -3948
rect 10761 -3914 12641 -3898
rect 10761 -3948 10777 -3914
rect 12625 -3948 12641 -3914
rect 10761 -3986 12641 -3948
rect 12699 -3914 14579 -3898
rect 12699 -3948 12715 -3914
rect 14563 -3948 14579 -3914
rect 12699 -3986 14579 -3948
rect 6885 -4324 8765 -4286
rect 6885 -4358 6901 -4324
rect 8749 -4358 8765 -4324
rect 6885 -4396 8765 -4358
rect 8823 -4324 10703 -4286
rect 8823 -4358 8839 -4324
rect 10687 -4358 10703 -4324
rect 8823 -4396 10703 -4358
rect 10761 -4324 12641 -4286
rect 10761 -4358 10777 -4324
rect 12625 -4358 12641 -4324
rect 10761 -4396 12641 -4358
rect 12699 -4324 14579 -4286
rect 12699 -4358 12715 -4324
rect 14563 -4358 14579 -4324
rect 12699 -4396 14579 -4358
rect 6885 -4734 8765 -4696
rect 6885 -4768 6901 -4734
rect 8749 -4768 8765 -4734
rect 6885 -4784 8765 -4768
rect 8823 -4734 10703 -4696
rect 8823 -4768 8839 -4734
rect 10687 -4768 10703 -4734
rect 8823 -4784 10703 -4768
rect 10761 -4734 12641 -4696
rect 10761 -4768 10777 -4734
rect 12625 -4768 12641 -4734
rect 10761 -4784 12641 -4768
rect 12699 -4734 14579 -4696
rect 12699 -4768 12715 -4734
rect 14563 -4768 14579 -4734
rect 12699 -4784 14579 -4768
<< polycont >>
rect 6891 4064 7239 4098
rect 7329 4064 7677 4098
rect 7767 4064 8115 4098
rect 8205 4064 8553 4098
rect 6891 936 7239 970
rect 7329 936 7677 970
rect 7767 936 8115 970
rect 8205 936 8553 970
rect 6891 87 7239 121
rect 7329 87 7677 121
rect 7767 87 8115 121
rect 8205 87 8553 121
rect 6891 -3041 7239 -3007
rect 7329 -3041 7677 -3007
rect 7767 -3041 8115 -3007
rect 8205 -3041 8553 -3007
rect 11720 -1467 12048 -1433
rect 12138 -1467 12466 -1433
rect 12556 -1467 12884 -1433
rect 12974 -1467 13302 -1433
rect 11720 -2995 12048 -2961
rect 12138 -2995 12466 -2961
rect 12556 -2995 12884 -2961
rect 12974 -2995 13302 -2961
rect 6901 -3948 8749 -3914
rect 8839 -3948 10687 -3914
rect 10777 -3948 12625 -3914
rect 12715 -3948 14563 -3914
rect 6901 -4358 8749 -4324
rect 8839 -4358 10687 -4324
rect 10777 -4358 12625 -4324
rect 12715 -4358 14563 -4324
rect 6901 -4768 8749 -4734
rect 8839 -4768 10687 -4734
rect 10777 -4768 12625 -4734
rect 12715 -4768 14563 -4734
<< xpolycontact >>
rect 14590 -1959 14660 -1527
rect 14590 -2559 14660 -2127
<< xpolyres >>
rect 14590 -2127 14660 -1959
<< locali >>
rect 6457 4501 9122 4514
rect 6457 890 6491 4501
rect 9083 4298 9122 4501
rect 6656 4280 8931 4298
rect 6656 890 6691 4280
rect 6875 4064 6891 4098
rect 7239 4064 7255 4098
rect 7313 4064 7329 4098
rect 7677 4064 7693 4098
rect 7751 4064 7767 4098
rect 8115 4064 8131 4098
rect 8189 4064 8205 4098
rect 8553 4064 8569 4098
rect 6829 4005 6863 4021
rect 6829 1013 6863 1029
rect 7267 4005 7301 4021
rect 7267 1013 7301 1029
rect 7705 4005 7739 4021
rect 7705 1013 7739 1029
rect 8143 4005 8177 4021
rect 8143 1013 8177 1029
rect 8581 4005 8615 4021
rect 8581 1013 8615 1029
rect 8806 3719 8931 4280
rect 8965 3719 9122 4298
rect 8806 1239 8871 3719
rect 9013 1239 9122 3719
rect 6875 936 6891 970
rect 7239 936 7255 970
rect 7313 936 7329 970
rect 7677 936 7693 970
rect 7751 936 7767 970
rect 8115 936 8131 970
rect 8189 936 8205 970
rect 8553 936 8569 970
rect 6457 72 6565 890
rect 6599 72 6691 890
rect 6875 87 6891 121
rect 7239 87 7255 121
rect 7313 87 7329 121
rect 7677 87 7693 121
rect 7751 87 7767 121
rect 8115 87 8131 121
rect 8189 87 8205 121
rect 8553 87 8569 121
rect 6457 -3104 6508 72
rect 6457 -3280 6507 -3104
rect 6656 -3123 6691 72
rect 6829 28 6863 44
rect 6829 -2964 6863 -2948
rect 7267 28 7301 44
rect 7267 -2964 7301 -2948
rect 7705 28 7739 44
rect 7705 -2964 7739 -2948
rect 8143 28 8177 44
rect 8143 -2964 8177 -2948
rect 8581 28 8615 44
rect 8581 -2964 8615 -2948
rect 8806 -514 8931 1239
rect 8965 -514 9122 1239
rect 8806 -2994 8887 -514
rect 9029 -925 9122 -514
rect 9029 -1012 13862 -925
rect 13819 -1013 13862 -1012
rect 9029 -1391 11291 -1304
rect 9029 -2994 9122 -1391
rect 6875 -3041 6891 -3007
rect 7239 -3041 7255 -3007
rect 7313 -3041 7329 -3007
rect 7677 -3041 7693 -3007
rect 7751 -3041 7767 -3007
rect 8115 -3041 8131 -3007
rect 8189 -3041 8205 -3007
rect 8553 -3041 8569 -3007
rect 8806 -3123 8931 -2994
rect 6656 -3137 8931 -3123
rect 8965 -3137 9122 -2994
rect 9072 -3261 9122 -3137
rect 6457 -3281 6620 -3280
rect 9072 -3281 9108 -3261
rect 6457 -3288 9108 -3281
rect 11246 -3294 11291 -1391
rect 11524 -1331 13542 -1304
rect 11524 -1365 11640 -1331
rect 13382 -1365 13542 -1331
rect 11524 -1391 13542 -1365
rect 11524 -1427 11588 -1391
rect 11524 -3001 11544 -1427
rect 11578 -3001 11588 -1427
rect 13428 -1427 13542 -1391
rect 11704 -1467 11720 -1433
rect 12048 -1467 12064 -1433
rect 12122 -1467 12138 -1433
rect 12466 -1467 12482 -1433
rect 12540 -1467 12556 -1433
rect 12884 -1467 12900 -1433
rect 12958 -1467 12974 -1433
rect 13302 -1467 13318 -1433
rect 11658 -1526 11692 -1510
rect 11658 -2918 11692 -2902
rect 12076 -1526 12110 -1510
rect 12076 -2918 12110 -2902
rect 12494 -1526 12528 -1510
rect 12494 -2918 12528 -2902
rect 12912 -1526 12946 -1510
rect 12912 -2918 12946 -2902
rect 13330 -1526 13364 -1510
rect 13330 -2918 13364 -2902
rect 11704 -2995 11720 -2961
rect 12048 -2995 12064 -2961
rect 12122 -2995 12138 -2961
rect 12466 -2995 12482 -2961
rect 12540 -2995 12556 -2961
rect 12884 -2995 12900 -2961
rect 12958 -2995 12974 -2961
rect 13302 -2995 13318 -2961
rect 11524 -3034 11588 -3001
rect 13428 -3001 13444 -1427
rect 13478 -2820 13542 -1427
rect 13829 -2820 13862 -1013
rect 13478 -3001 13862 -2820
rect 13428 -3034 13862 -3001
rect 11524 -3054 13862 -3034
rect 14372 -1377 14889 -1350
rect 14372 -2526 14406 -1377
rect 14492 -1381 14889 -1377
rect 14492 -1397 14769 -1381
rect 14492 -1431 14556 -1397
rect 14694 -1431 14769 -1397
rect 14492 -1436 14769 -1431
rect 14492 -1493 14529 -1436
rect 14372 -2593 14460 -2526
rect 14494 -2593 14529 -1493
rect 14732 -1493 14769 -1436
rect 14372 -2622 14529 -2593
rect 11524 -3060 13866 -3054
rect 11246 -3296 11376 -3294
rect 13439 -3296 13866 -3060
rect 11246 -3310 13866 -3296
rect 14372 -3582 14389 -2622
rect 6553 -3619 14389 -3582
rect 6553 -5119 6563 -3619
rect 6710 -3622 14389 -3619
rect 14505 -2632 14529 -2622
rect 14732 -2593 14756 -1493
rect 14732 -2632 14769 -2593
rect 14505 -2655 14769 -2632
rect 14505 -2689 14556 -2655
rect 14694 -2689 14769 -2655
rect 14505 -2690 14769 -2689
rect 14848 -2690 14889 -1381
rect 14505 -2718 14889 -2690
rect 14505 -3582 14529 -2718
rect 14505 -3622 14960 -3582
rect 14846 -3656 14960 -3622
rect 14505 -3682 14960 -3656
rect 6710 -3743 14389 -3731
rect 14505 -3743 14872 -3682
rect 6710 -3769 14872 -3743
rect 6710 -4847 6731 -3769
rect 6885 -3948 6901 -3914
rect 8749 -3948 8765 -3914
rect 8823 -3948 8839 -3914
rect 10687 -3948 10703 -3914
rect 10761 -3948 10777 -3914
rect 12625 -3948 12641 -3914
rect 12699 -3948 12715 -3914
rect 14563 -3948 14579 -3914
rect 6839 -3998 6873 -3982
rect 6839 -4290 6873 -4274
rect 8777 -3998 8811 -3982
rect 8777 -4290 8811 -4274
rect 10715 -3998 10749 -3982
rect 10715 -4290 10749 -4274
rect 12653 -3998 12687 -3982
rect 12653 -4290 12687 -4274
rect 14591 -3998 14625 -3982
rect 14591 -4290 14625 -4274
rect 6885 -4358 6901 -4324
rect 8749 -4358 8765 -4324
rect 8823 -4358 8839 -4324
rect 10687 -4358 10703 -4324
rect 10761 -4358 10777 -4324
rect 12625 -4358 12641 -4324
rect 12699 -4358 12715 -4324
rect 14563 -4358 14579 -4324
rect 6839 -4408 6873 -4392
rect 6839 -4700 6873 -4684
rect 8777 -4408 8811 -4392
rect 8777 -4700 8811 -4684
rect 10715 -4408 10749 -4392
rect 10715 -4700 10749 -4684
rect 12653 -4408 12687 -4392
rect 12653 -4700 12687 -4684
rect 14591 -4408 14625 -4392
rect 14591 -4700 14625 -4684
rect 6885 -4768 6901 -4734
rect 8749 -4768 8765 -4734
rect 8823 -4768 8839 -4734
rect 10687 -4768 10703 -4734
rect 10761 -4768 10777 -4734
rect 12625 -4768 12641 -4734
rect 12699 -4768 12715 -4734
rect 14563 -4768 14579 -4734
rect 14791 -4847 14872 -3769
rect 6710 -4905 14872 -4847
rect 14906 -4905 14960 -3682
rect 6710 -4921 14960 -4905
rect 6804 -4922 14960 -4921
rect 14482 -4931 14960 -4922
rect 14846 -4965 14960 -4931
rect 14482 -5119 14960 -4965
rect 6553 -5136 14960 -5119
rect 6562 -5137 14960 -5136
<< viali >>
rect 6491 4431 9083 4501
rect 6491 4397 6625 4431
rect 6625 4397 8905 4431
rect 8905 4397 9083 4431
rect 6491 4371 9083 4397
rect 6491 890 6565 4371
rect 6565 890 6599 4371
rect 6599 4298 8931 4371
rect 8931 4298 8965 4371
rect 8965 4298 9083 4371
rect 6599 890 6656 4298
rect 6891 4064 7239 4098
rect 7329 4064 7677 4098
rect 7767 4064 8115 4098
rect 8205 4064 8553 4098
rect 6829 1029 6863 4005
rect 7267 1029 7301 4005
rect 7705 1029 7739 4005
rect 8143 1029 8177 4005
rect 8581 1029 8615 4005
rect 8871 1239 8931 3719
rect 8931 1239 8965 3719
rect 8965 1239 9013 3719
rect 6891 936 7239 970
rect 7329 936 7677 970
rect 7767 936 8115 970
rect 8205 936 8553 970
rect 6891 87 7239 121
rect 7329 87 7677 121
rect 7767 87 8115 121
rect 8205 87 8553 121
rect 6508 -3104 6565 72
rect 6507 -3164 6565 -3104
rect 6565 -3164 6599 72
rect 6599 -3137 6656 72
rect 6829 -2948 6863 28
rect 7267 -2948 7301 28
rect 7705 -2948 7739 28
rect 8143 -2948 8177 28
rect 8581 -2948 8615 28
rect 8887 -2994 8931 -514
rect 8931 -2994 8965 -514
rect 8965 -1012 9029 -514
rect 8965 -1013 13819 -1012
rect 8965 -1304 13829 -1013
rect 8965 -2994 9029 -1304
rect 6891 -3041 7239 -3007
rect 7329 -3041 7677 -3007
rect 7767 -3041 8115 -3007
rect 8205 -3041 8553 -3007
rect 6599 -3164 8931 -3137
rect 8931 -3164 8965 -3137
rect 8965 -3164 9072 -3137
rect 6507 -3190 9072 -3164
rect 6507 -3224 6625 -3190
rect 6625 -3224 8905 -3190
rect 8905 -3224 9072 -3190
rect 6507 -3280 9072 -3224
rect 6620 -3281 9072 -3280
rect 11291 -3060 11524 -1304
rect 11720 -1467 12048 -1433
rect 12138 -1467 12466 -1433
rect 12556 -1467 12884 -1433
rect 12974 -1467 13302 -1433
rect 11658 -2902 11692 -1526
rect 12076 -2902 12110 -1526
rect 12494 -2902 12528 -1526
rect 12912 -2902 12946 -1526
rect 13330 -2902 13364 -1526
rect 11720 -2995 12048 -2961
rect 12138 -2995 12466 -2961
rect 12556 -2995 12884 -2961
rect 12974 -2995 13302 -2961
rect 13542 -2820 13829 -1304
rect 14406 -1493 14492 -1377
rect 14406 -2526 14460 -1493
rect 14460 -2526 14492 -1493
rect 14769 -1493 14848 -1381
rect 14606 -1942 14644 -1545
rect 14606 -2541 14644 -2144
rect 11291 -3063 13439 -3060
rect 11291 -3097 11640 -3063
rect 11640 -3097 13382 -3063
rect 13382 -3097 13439 -3063
rect 11291 -3294 13439 -3097
rect 11376 -3296 13439 -3294
rect 6563 -3622 6710 -3619
rect 14389 -3622 14505 -2622
rect 14769 -2593 14790 -1493
rect 14790 -2593 14848 -1493
rect 14769 -2690 14848 -2593
rect 6563 -3656 6677 -3622
rect 6677 -3627 6710 -3622
rect 6677 -3628 6839 -3627
rect 14389 -3628 14505 -3622
rect 6677 -3656 14505 -3628
rect 6563 -3682 14505 -3656
rect 6563 -4905 6617 -3682
rect 6617 -4905 6651 -3682
rect 6651 -3731 14505 -3682
rect 6651 -4905 6710 -3731
rect 14389 -3743 14505 -3731
rect 6901 -3948 8749 -3914
rect 8839 -3948 10687 -3914
rect 10777 -3948 12625 -3914
rect 12715 -3948 14563 -3914
rect 6839 -4274 6873 -3998
rect 8777 -4274 8811 -3998
rect 10715 -4274 10749 -3998
rect 12653 -4274 12687 -3998
rect 14591 -4274 14625 -3998
rect 6901 -4358 8749 -4324
rect 8839 -4358 10687 -4324
rect 10777 -4358 12625 -4324
rect 12715 -4358 14563 -4324
rect 6839 -4684 6873 -4408
rect 8777 -4684 8811 -4408
rect 10715 -4684 10749 -4408
rect 12653 -4684 12687 -4408
rect 14591 -4684 14625 -4408
rect 6901 -4768 8749 -4734
rect 8839 -4768 10687 -4734
rect 10777 -4768 12625 -4734
rect 12715 -4768 14563 -4734
rect 6563 -4921 6710 -4905
rect 6563 -4922 6804 -4921
rect 6563 -4931 14482 -4922
rect 6563 -4965 6677 -4931
rect 6677 -4965 14482 -4931
rect 6563 -5119 14482 -4965
<< metal1 >>
rect 6479 4501 9095 4507
rect 6479 4292 6491 4501
rect 9083 4298 9095 4501
rect 6481 890 6491 4292
rect 6656 4292 9095 4298
rect 6656 890 6666 4292
rect 6879 4098 7251 4104
rect 6879 4064 6891 4098
rect 7239 4064 7251 4098
rect 6879 4058 7251 4064
rect 7317 4098 7689 4104
rect 7317 4064 7329 4098
rect 7677 4064 7689 4098
rect 7317 4058 7689 4064
rect 7755 4098 8127 4104
rect 7755 4064 7767 4098
rect 8115 4064 8127 4098
rect 7755 4058 8127 4064
rect 8193 4098 8565 4104
rect 8193 4064 8205 4098
rect 8553 4064 8565 4098
rect 8193 4058 8565 4064
rect 6823 4005 6869 4017
rect 6823 2029 6829 4005
rect 6863 2029 6869 4005
rect 6803 1029 6813 2029
rect 6877 1029 6887 2029
rect 6823 1017 6869 1029
rect 6951 979 7156 4058
rect 7261 4005 7307 4017
rect 7238 3405 7248 4005
rect 7320 3405 7330 4005
rect 7261 1029 7267 3405
rect 7301 1029 7307 3405
rect 7261 1017 7307 1029
rect 7404 979 7609 4058
rect 7699 4005 7745 4017
rect 7699 3266 7705 4005
rect 7739 3266 7745 4005
rect 7680 2266 7690 3266
rect 7754 2266 7764 3266
rect 7699 1029 7705 2266
rect 7739 1029 7745 2266
rect 7699 1017 7745 1029
rect 7840 979 8045 4058
rect 8137 4005 8183 4017
rect 8114 3405 8124 4005
rect 8196 3405 8206 4005
rect 8137 1029 8143 3405
rect 8177 1029 8183 3405
rect 8137 1017 8183 1029
rect 8280 979 8485 4058
rect 8575 4005 8621 4017
rect 8575 2029 8581 4005
rect 8615 2029 8621 4005
rect 8865 3719 9019 3731
rect 8556 1029 8566 2029
rect 8630 1029 8640 2029
rect 8865 1239 8871 3719
rect 9013 1239 9019 3719
rect 8865 1227 9019 1239
rect 8575 1017 8621 1029
rect 6881 976 6891 979
rect 6879 930 6891 976
rect 7171 976 7181 979
rect 7319 976 7329 979
rect 7171 970 7251 976
rect 7239 936 7251 970
rect 6881 927 6891 930
rect 7171 930 7251 936
rect 7317 930 7329 976
rect 7609 976 7619 979
rect 7757 976 7767 979
rect 7609 970 7689 976
rect 7677 936 7689 970
rect 7171 927 7181 930
rect 7319 927 7329 930
rect 7609 930 7689 936
rect 7755 930 7767 976
rect 8047 976 8057 979
rect 8195 976 8205 979
rect 8047 970 8127 976
rect 8115 936 8127 970
rect 7609 927 7619 930
rect 7757 927 7767 930
rect 8047 930 8127 936
rect 8193 930 8205 976
rect 8485 976 8495 979
rect 8485 970 8565 976
rect 8553 936 8565 970
rect 8047 927 8057 930
rect 8195 927 8205 930
rect 8485 930 8565 936
rect 8485 927 8495 930
rect 6485 878 6662 890
rect 6296 634 6891 734
rect 6991 634 7577 734
rect 7677 634 8015 734
rect 8115 634 8205 734
rect 8305 634 10030 734
rect 10312 634 10322 734
rect 6296 325 7139 425
rect 7239 325 7329 425
rect 7429 325 7767 425
rect 7867 325 8453 425
rect 8553 325 8710 425
rect 6949 127 6959 130
rect 6879 121 6959 127
rect 7239 127 7249 130
rect 7387 127 7397 130
rect 6879 87 6891 121
rect 6502 72 6662 84
rect 6879 81 6959 87
rect 6949 78 6959 81
rect 7239 81 7251 127
rect 7317 121 7397 127
rect 7677 127 7687 130
rect 7825 127 7835 130
rect 7317 87 7329 121
rect 7317 81 7397 87
rect 7239 78 7249 81
rect 7387 78 7397 81
rect 7677 81 7689 127
rect 7755 121 7835 127
rect 8115 127 8125 130
rect 8263 127 8273 130
rect 7755 87 7767 121
rect 7755 81 7835 87
rect 7677 78 7687 81
rect 7825 78 7835 81
rect 8115 81 8127 127
rect 8193 121 8273 127
rect 8553 127 8563 130
rect 8193 87 8205 121
rect 8193 81 8273 87
rect 8115 78 8125 81
rect 8263 78 8273 81
rect 8553 81 8565 127
rect 8553 78 8563 81
rect 6498 -3104 6508 72
rect 6497 -3280 6507 -3104
rect 6656 -3131 6666 72
rect 6823 28 6869 40
rect 6804 -972 6814 28
rect 6878 -972 6888 28
rect 6823 -2948 6829 -972
rect 6863 -2948 6869 -972
rect 6823 -2960 6869 -2948
rect 6955 -3001 7160 78
rect 7261 28 7307 40
rect 7261 -2348 7267 28
rect 7301 -2348 7307 28
rect 7238 -2948 7248 -2348
rect 7320 -2948 7330 -2348
rect 7261 -2960 7307 -2948
rect 7408 -3001 7613 78
rect 7699 28 7745 40
rect 7699 -1132 7705 28
rect 7739 -1132 7745 28
rect 7680 -2132 7690 -1132
rect 7754 -2132 7764 -1132
rect 7699 -2948 7705 -2132
rect 7739 -2948 7745 -2132
rect 7699 -2960 7745 -2948
rect 7844 -3001 8049 78
rect 8137 28 8183 40
rect 8137 -2348 8143 28
rect 8177 -2348 8183 28
rect 8113 -2948 8123 -2348
rect 8195 -2948 8205 -2348
rect 8137 -2960 8183 -2948
rect 8276 -3001 8481 78
rect 8575 28 8621 40
rect 8556 -972 8566 28
rect 8630 -972 8640 28
rect 8881 -514 9035 -502
rect 8575 -2948 8581 -972
rect 8615 -2948 8621 -972
rect 8575 -2960 8621 -2948
rect 8881 -2994 8887 -514
rect 9029 -1006 9035 -514
rect 13536 -1006 13835 -1001
rect 9029 -1012 13835 -1006
rect 13819 -1013 13835 -1012
rect 9029 -1310 11291 -1304
rect 9029 -2994 9035 -1310
rect 6879 -3007 7251 -3001
rect 6879 -3041 6891 -3007
rect 7239 -3041 7251 -3007
rect 6879 -3047 7251 -3041
rect 7317 -3007 7689 -3001
rect 7317 -3041 7329 -3007
rect 7677 -3041 7689 -3007
rect 7317 -3047 7689 -3041
rect 7755 -3007 8127 -3001
rect 7755 -3041 7767 -3007
rect 8115 -3041 8127 -3007
rect 7755 -3047 8127 -3041
rect 8193 -3007 8565 -3001
rect 8881 -3006 9035 -2994
rect 8193 -3041 8205 -3007
rect 8553 -3041 8565 -3007
rect 8193 -3047 8565 -3041
rect 6656 -3137 9084 -3131
rect 6501 -3281 6620 -3280
rect 9072 -3281 9084 -3137
rect 6501 -3287 9084 -3281
rect 6501 -3292 6662 -3287
rect 11285 -3294 11291 -1310
rect 11524 -1310 13542 -1304
rect 11524 -3054 11530 -1310
rect 11708 -1433 12060 -1427
rect 11708 -1467 11720 -1433
rect 12048 -1467 12060 -1433
rect 11708 -1473 12060 -1467
rect 12126 -1433 12478 -1427
rect 12126 -1467 12138 -1433
rect 12466 -1467 12478 -1433
rect 12126 -1473 12478 -1467
rect 12544 -1433 12896 -1427
rect 12544 -1467 12556 -1433
rect 12884 -1467 12896 -1433
rect 12544 -1473 12896 -1467
rect 12962 -1433 13314 -1427
rect 12962 -1467 12974 -1433
rect 13302 -1467 13314 -1433
rect 12962 -1473 13314 -1467
rect 11652 -1526 11698 -1514
rect 11639 -2526 11649 -1526
rect 11701 -2526 11711 -1526
rect 11652 -2902 11658 -2526
rect 11692 -2902 11698 -2526
rect 11652 -2914 11698 -2902
rect 11776 -2955 11977 -1473
rect 12070 -1526 12116 -1514
rect 12070 -1902 12076 -1526
rect 12110 -1902 12116 -1526
rect 12057 -2902 12067 -1902
rect 12119 -2902 12129 -1902
rect 12070 -2914 12116 -2902
rect 12195 -2955 12396 -1473
rect 12488 -1526 12534 -1514
rect 12475 -2526 12485 -1526
rect 12537 -2526 12547 -1526
rect 12488 -2902 12494 -2526
rect 12528 -2902 12534 -2526
rect 12488 -2914 12534 -2902
rect 12618 -2955 12819 -1473
rect 12906 -1526 12952 -1514
rect 12906 -1902 12912 -1526
rect 12946 -1902 12952 -1526
rect 12893 -2902 12903 -1902
rect 12955 -2902 12965 -1902
rect 12906 -2914 12952 -2902
rect 13024 -2955 13225 -1473
rect 13324 -1526 13370 -1514
rect 13311 -2526 13321 -1526
rect 13373 -2526 13383 -1526
rect 13324 -2902 13330 -2526
rect 13364 -2902 13370 -2526
rect 13532 -2820 13542 -1310
rect 13829 -2820 13839 -1013
rect 14400 -1377 14498 -1365
rect 14396 -2526 14406 -1377
rect 14492 -2526 14502 -1377
rect 14763 -1381 14854 -1369
rect 14600 -1545 14650 -1533
rect 14583 -1665 14593 -1545
rect 14657 -1665 14667 -1545
rect 14600 -1942 14606 -1665
rect 14644 -1942 14650 -1665
rect 14600 -1954 14650 -1942
rect 14600 -2144 14650 -2132
rect 14600 -2421 14606 -2144
rect 14644 -2421 14650 -2144
rect 14400 -2538 14498 -2526
rect 14582 -2541 14592 -2421
rect 14656 -2541 14666 -2421
rect 14600 -2553 14650 -2541
rect 14383 -2622 14511 -2610
rect 13536 -2832 13835 -2820
rect 13324 -2914 13370 -2902
rect 13519 -2955 13529 -2946
rect 11708 -2961 13529 -2955
rect 11708 -2995 11720 -2961
rect 12048 -2995 12138 -2961
rect 12466 -2995 12556 -2961
rect 12884 -2995 12974 -2961
rect 13302 -2995 13529 -2961
rect 11708 -3001 13529 -2995
rect 13519 -3005 13529 -3001
rect 13653 -3005 13663 -2946
rect 11524 -3060 13451 -3054
rect 11285 -3296 11376 -3294
rect 13439 -3296 13451 -3060
rect 11285 -3302 13451 -3296
rect 11285 -3306 11530 -3302
rect 6557 -3619 6716 -3607
rect 6553 -4915 6563 -3619
rect 6710 -3621 6720 -3619
rect 6710 -3622 6851 -3621
rect 14383 -3622 14389 -2622
rect 6710 -3627 14389 -3622
rect 6839 -3628 14389 -3627
rect 6551 -5119 6563 -4915
rect 6710 -3737 14389 -3731
rect 6710 -4915 6720 -3737
rect 14383 -3743 14389 -3737
rect 14505 -3743 14511 -2622
rect 14759 -2690 14769 -1381
rect 14848 -2690 14858 -1381
rect 14763 -2702 14854 -2690
rect 14383 -3755 14511 -3743
rect 6889 -3914 8761 -3908
rect 6889 -3948 6901 -3914
rect 8749 -3948 8761 -3914
rect 6889 -3954 8761 -3948
rect 8827 -3914 12637 -3908
rect 8827 -3948 8839 -3914
rect 10687 -3948 10777 -3914
rect 12625 -3948 12637 -3914
rect 8827 -3954 12637 -3948
rect 12703 -3914 14575 -3908
rect 12703 -3948 12715 -3914
rect 14563 -3948 14575 -3914
rect 12703 -3954 14575 -3948
rect 6833 -3998 6879 -3986
rect 6814 -4098 6824 -3998
rect 6888 -4098 6898 -3998
rect 6833 -4274 6839 -4098
rect 6873 -4274 6879 -4098
rect 6833 -4286 6879 -4274
rect 7109 -4318 8528 -3954
rect 8771 -3998 8817 -3986
rect 8758 -4098 8768 -3998
rect 8820 -4098 8830 -3998
rect 8771 -4274 8777 -4098
rect 8811 -4274 8817 -4098
rect 8771 -4286 8817 -4274
rect 9143 -4318 10562 -3954
rect 10709 -3998 10755 -3954
rect 10709 -4174 10715 -3998
rect 10749 -4174 10755 -3998
rect 10690 -4274 10700 -4174
rect 10764 -4274 10774 -4174
rect 10709 -4286 10755 -4274
rect 10972 -4318 12391 -3954
rect 12647 -3998 12693 -3986
rect 12634 -4098 12644 -3998
rect 12696 -4098 12706 -3998
rect 12647 -4274 12653 -4098
rect 12687 -4274 12693 -4098
rect 12647 -4286 12693 -4274
rect 12942 -4318 14361 -3954
rect 14585 -3998 14631 -3986
rect 14566 -4098 14576 -3998
rect 14640 -4098 14650 -3998
rect 14585 -4274 14591 -4098
rect 14625 -4274 14631 -4098
rect 14585 -4286 14631 -4274
rect 6889 -4324 14575 -4318
rect 6889 -4358 6901 -4324
rect 8749 -4358 8839 -4324
rect 10687 -4358 10777 -4324
rect 12625 -4358 12715 -4324
rect 14563 -4358 14575 -4324
rect 6889 -4364 14575 -4358
rect 6833 -4408 6879 -4396
rect 6833 -4584 6839 -4408
rect 6873 -4584 6879 -4408
rect 6814 -4684 6824 -4584
rect 6888 -4684 6898 -4584
rect 6833 -4728 6879 -4684
rect 7113 -4728 8532 -4364
rect 8771 -4408 8817 -4396
rect 8771 -4584 8777 -4408
rect 8811 -4584 8817 -4408
rect 8758 -4684 8768 -4584
rect 8820 -4684 8830 -4584
rect 8771 -4696 8817 -4684
rect 9139 -4728 10558 -4364
rect 10709 -4408 10755 -4396
rect 10690 -4508 10700 -4408
rect 10764 -4508 10774 -4408
rect 10709 -4684 10715 -4508
rect 10749 -4684 10755 -4508
rect 10709 -4696 10755 -4684
rect 10972 -4728 12391 -4364
rect 12647 -4408 12693 -4396
rect 12647 -4584 12653 -4408
rect 12687 -4584 12693 -4408
rect 12634 -4684 12644 -4584
rect 12696 -4684 12706 -4584
rect 12647 -4696 12693 -4684
rect 12942 -4728 14361 -4364
rect 14585 -4408 14631 -4396
rect 14585 -4584 14591 -4408
rect 14625 -4584 14631 -4408
rect 14566 -4684 14576 -4584
rect 14640 -4684 14650 -4584
rect 14585 -4728 14631 -4684
rect 6833 -4734 8761 -4728
rect 6833 -4768 6901 -4734
rect 8749 -4768 8761 -4734
rect 6833 -4774 8761 -4768
rect 8827 -4734 10699 -4728
rect 8827 -4768 8839 -4734
rect 10687 -4768 10699 -4734
rect 8827 -4774 10699 -4768
rect 10765 -4734 12637 -4728
rect 10765 -4768 10777 -4734
rect 12625 -4768 12637 -4734
rect 10765 -4774 12637 -4768
rect 12703 -4734 14631 -4728
rect 12703 -4768 12715 -4734
rect 14563 -4768 14631 -4734
rect 12703 -4774 14631 -4768
rect 6710 -4916 6816 -4915
rect 6710 -4921 14494 -4916
rect 6804 -4922 14494 -4921
rect 14482 -5119 14494 -4922
rect 6551 -5125 14494 -5119
<< via1 >>
rect 6491 4298 9083 4501
rect 6491 890 6656 4298
rect 6813 1029 6829 2029
rect 6829 1029 6863 2029
rect 6863 1029 6877 2029
rect 7248 3405 7267 4005
rect 7267 3405 7301 4005
rect 7301 3405 7320 4005
rect 7690 2266 7705 3266
rect 7705 2266 7739 3266
rect 7739 2266 7754 3266
rect 8124 3405 8143 4005
rect 8143 3405 8177 4005
rect 8177 3405 8196 4005
rect 8566 1029 8581 2029
rect 8581 1029 8615 2029
rect 8615 1029 8630 2029
rect 6891 970 7171 979
rect 6891 936 7171 970
rect 6891 927 7171 936
rect 7329 970 7609 979
rect 7329 936 7609 970
rect 7329 927 7609 936
rect 7767 970 8047 979
rect 7767 936 8047 970
rect 7767 927 8047 936
rect 8205 970 8485 979
rect 8205 936 8485 970
rect 8205 927 8485 936
rect 6891 634 6991 734
rect 7577 634 7677 734
rect 8015 634 8115 734
rect 8205 634 8305 734
rect 10030 634 10312 734
rect 7139 325 7239 425
rect 7329 325 7429 425
rect 7767 325 7867 425
rect 8453 325 8553 425
rect 6959 121 7239 130
rect 6959 87 7239 121
rect 6959 78 7239 87
rect 7397 121 7677 130
rect 7397 87 7677 121
rect 7397 78 7677 87
rect 7835 121 8115 130
rect 7835 87 8115 121
rect 7835 78 8115 87
rect 8273 121 8553 130
rect 8273 87 8553 121
rect 8273 78 8553 87
rect 6508 -3104 6656 72
rect 6507 -3137 6656 -3104
rect 6814 -972 6829 28
rect 6829 -972 6863 28
rect 6863 -972 6878 28
rect 7248 -2948 7267 -2348
rect 7267 -2948 7301 -2348
rect 7301 -2948 7320 -2348
rect 7690 -2132 7705 -1132
rect 7705 -2132 7739 -1132
rect 7739 -2132 7754 -1132
rect 8123 -2948 8143 -2348
rect 8143 -2948 8177 -2348
rect 8177 -2948 8195 -2348
rect 8566 -972 8581 28
rect 8581 -972 8615 28
rect 8615 -972 8630 28
rect 10166 -1304 13829 -1013
rect 6507 -3280 9072 -3137
rect 6620 -3281 9072 -3280
rect 11649 -2526 11658 -1526
rect 11658 -2526 11692 -1526
rect 11692 -2526 11701 -1526
rect 12067 -2902 12076 -1902
rect 12076 -2902 12110 -1902
rect 12110 -2902 12119 -1902
rect 12485 -2526 12494 -1526
rect 12494 -2526 12528 -1526
rect 12528 -2526 12537 -1526
rect 12903 -2902 12912 -1902
rect 12912 -2902 12946 -1902
rect 12946 -2902 12955 -1902
rect 13321 -2526 13330 -1526
rect 13330 -2526 13364 -1526
rect 13364 -2526 13373 -1526
rect 13542 -2820 13829 -1304
rect 14406 -2526 14492 -1377
rect 14593 -1665 14606 -1545
rect 14606 -1665 14644 -1545
rect 14644 -1665 14657 -1545
rect 14592 -2541 14606 -2421
rect 14606 -2541 14644 -2421
rect 14644 -2541 14656 -2421
rect 13529 -3005 13653 -2946
rect 11376 -3296 13439 -3060
rect 6563 -3627 6710 -3619
rect 6563 -3628 6839 -3627
rect 6563 -3731 14454 -3628
rect 6563 -4921 6710 -3731
rect 14769 -2690 14848 -1381
rect 6824 -4098 6839 -3998
rect 6839 -4098 6873 -3998
rect 6873 -4098 6888 -3998
rect 8768 -4098 8777 -3998
rect 8777 -4098 8811 -3998
rect 8811 -4098 8820 -3998
rect 10700 -4274 10715 -4174
rect 10715 -4274 10749 -4174
rect 10749 -4274 10764 -4174
rect 12644 -4098 12653 -3998
rect 12653 -4098 12687 -3998
rect 12687 -4098 12696 -3998
rect 14576 -4098 14591 -3998
rect 14591 -4098 14625 -3998
rect 14625 -4098 14640 -3998
rect 6824 -4684 6839 -4584
rect 6839 -4684 6873 -4584
rect 6873 -4684 6888 -4584
rect 8768 -4684 8777 -4584
rect 8777 -4684 8811 -4584
rect 8811 -4684 8820 -4584
rect 10700 -4508 10715 -4408
rect 10715 -4508 10749 -4408
rect 10749 -4508 10764 -4408
rect 12644 -4684 12653 -4584
rect 12653 -4684 12687 -4584
rect 12687 -4684 12696 -4584
rect 14576 -4684 14591 -4584
rect 14591 -4684 14625 -4584
rect 14625 -4684 14640 -4584
rect 6563 -4922 6804 -4921
rect 6563 -5119 14482 -4922
<< metal2 >>
rect 6402 4501 9083 4511
rect 6402 4287 6491 4501
rect 6656 4288 9083 4298
rect 7248 4005 9929 4015
rect 7320 3915 8124 4005
rect 7248 3395 7320 3405
rect 8196 3915 9929 4005
rect 8124 3395 8196 3405
rect 7690 3266 7754 3276
rect 7690 2256 7754 2266
rect 6813 2029 6877 2039
rect 6813 1019 6877 1029
rect 8566 2029 8630 2039
rect 8566 1019 8630 1029
rect 6491 880 6656 890
rect 6891 979 7171 989
rect 6891 917 7171 927
rect 7329 979 7609 989
rect 7329 917 7609 927
rect 7767 979 8047 989
rect 7767 917 8047 927
rect 8205 979 8485 989
rect 8205 917 8485 927
rect 6891 734 6991 917
rect 6891 624 6991 634
rect 7139 425 7239 435
rect 7139 140 7239 325
rect 7329 425 7429 917
rect 7329 315 7429 325
rect 7577 734 7677 744
rect 7577 140 7677 634
rect 7767 425 7867 917
rect 7767 315 7867 325
rect 8015 734 8115 744
rect 8015 140 8115 634
rect 8205 734 8305 917
rect 8205 624 8305 634
rect 8453 425 8553 435
rect 8453 140 8553 325
rect 6959 130 7239 140
rect 6508 72 6656 82
rect 6507 -3104 6508 -3094
rect 6959 68 7239 78
rect 7397 130 7677 140
rect 7397 68 7677 78
rect 7835 130 8115 140
rect 7835 68 8115 78
rect 8273 130 8553 140
rect 8273 68 8553 78
rect 6814 28 6878 38
rect 6814 -982 6878 -972
rect 8566 28 8630 38
rect 8566 -982 8630 -972
rect 7690 -1132 7754 -1122
rect 7690 -2142 7754 -2132
rect 9829 -1516 9929 3915
rect 10020 734 10312 744
rect 10020 624 10312 634
rect 10166 -1013 13829 -1003
rect 10166 -1314 13542 -1304
rect 9829 -1526 13373 -1516
rect 9829 -1616 11649 -1526
rect 7248 -2338 8648 -2337
rect 9829 -2338 9929 -1616
rect 7248 -2348 9929 -2338
rect 7320 -2437 8123 -2348
rect 7248 -2958 7320 -2948
rect 8195 -2437 9929 -2348
rect 8520 -2438 9929 -2437
rect 11701 -1616 12485 -1526
rect 11649 -2536 11701 -2526
rect 12067 -1902 12119 -1892
rect 8123 -2958 8195 -2948
rect 12537 -1616 13321 -1526
rect 12485 -2536 12537 -2526
rect 12903 -1902 12955 -1892
rect 12067 -3050 12119 -2902
rect 13321 -2536 13373 -2526
rect 14406 -1377 14492 -1367
rect 14769 -1381 14848 -1371
rect 14593 -1545 14657 -1535
rect 14593 -1675 14657 -1665
rect 14406 -2536 14492 -2526
rect 14592 -2421 14656 -2411
rect 14592 -2551 14656 -2541
rect 14769 -2700 14848 -2690
rect 13542 -2830 13829 -2820
rect 12903 -3050 12955 -2902
rect 13529 -2946 15141 -2936
rect 13653 -3005 15141 -2946
rect 13529 -3015 15141 -3005
rect 11376 -3060 13439 -3050
rect 6656 -3137 9072 -3127
rect 6507 -3281 6620 -3280
rect 6507 -3290 9072 -3281
rect 6620 -3291 9072 -3290
rect 11376 -3306 13439 -3296
rect 6563 -3617 6710 -3609
rect 6563 -3618 6839 -3617
rect 6563 -3619 14454 -3618
rect 6710 -3627 14454 -3619
rect 6839 -3628 14454 -3627
rect 6497 -5119 6563 -4911
rect 6710 -3741 14454 -3731
rect 6824 -3998 6888 -3988
rect 6824 -4108 6888 -4098
rect 8768 -3998 8820 -3741
rect 8768 -4108 8820 -4098
rect 12644 -3998 12696 -3741
rect 12644 -4108 12696 -4098
rect 14576 -3998 14640 -3988
rect 14576 -4108 14640 -4098
rect 10700 -4174 10764 -4164
rect 10700 -4284 10764 -4274
rect 10700 -4408 10764 -4398
rect 10700 -4518 10764 -4508
rect 6824 -4584 6888 -4574
rect 6824 -4694 6888 -4684
rect 8768 -4584 8820 -4574
rect 6710 -4912 6804 -4911
rect 8768 -4912 8820 -4684
rect 12644 -4584 12696 -4574
rect 12644 -4912 12696 -4684
rect 14576 -4584 14640 -4574
rect 14576 -4694 14640 -4684
rect 6710 -4921 14482 -4912
rect 6804 -4922 14482 -4921
rect 15062 -5083 15141 -3015
rect 6497 -5129 14482 -5119
<< via2 >>
rect 7690 2266 7754 3266
rect 6813 1029 6877 2029
rect 8566 1029 8630 2029
rect 6814 -972 6878 28
rect 8566 -972 8630 28
rect 7690 -2132 7754 -1132
rect 10020 634 10030 734
rect 10030 634 10312 734
rect 14593 -1665 14657 -1545
rect 14592 -2541 14656 -2421
rect 6824 -4098 6888 -3998
rect 14576 -4098 14640 -3998
rect 10700 -4274 10764 -4174
rect 10700 -4508 10764 -4408
rect 6824 -4684 6888 -4584
rect 14576 -4684 14640 -4584
<< metal3 >>
rect 11255 4467 15627 4495
rect 7680 3266 7764 3271
rect 7680 2266 7690 3266
rect 7754 2352 7764 3266
rect 7754 2266 8872 2352
rect 7680 2261 8872 2266
rect 7694 2252 8872 2261
rect 6803 2029 6887 2034
rect 6803 1029 6813 2029
rect 6877 1029 6887 2029
rect 6803 1024 6887 1029
rect 8556 2029 8640 2034
rect 8556 1029 8566 2029
rect 8630 1029 8640 2029
rect 8556 1024 8640 1029
rect 8772 36 8872 2252
rect 11255 739 15543 4467
rect 10010 734 15543 739
rect 10010 634 10020 734
rect 10312 634 15543 734
rect 10010 629 15543 634
rect 11255 443 15543 629
rect 15607 443 15627 4467
rect 11255 415 15627 443
rect 8772 33 8963 36
rect 6804 28 8963 33
rect 6804 -972 6814 28
rect 6878 -67 8566 28
rect 6878 -972 6888 -67
rect 6804 -977 6888 -972
rect 8556 -972 8566 -67
rect 8630 -67 8963 28
rect 8630 -972 8640 -67
rect 8556 -977 8640 -972
rect 7680 -1132 7764 -1127
rect 7680 -2132 7690 -1132
rect 7754 -2132 7764 -1132
rect 7680 -2137 7764 -2132
rect 6807 -3998 6905 -3993
rect 6807 -4098 6824 -3998
rect 6888 -4098 6905 -3998
rect 6807 -4103 6905 -4098
rect 8853 -4169 8963 -67
rect 14583 -1545 14667 -1540
rect 14583 -1665 14593 -1545
rect 14657 -1665 14667 -1545
rect 14583 -1670 14667 -1665
rect 14582 -2421 14666 -2416
rect 14582 -2541 14592 -2421
rect 14656 -2541 14666 -2421
rect 14582 -2546 14666 -2541
rect 14538 -3998 14666 -3993
rect 14538 -4098 14576 -3998
rect 14640 -4098 14666 -3998
rect 14538 -4103 14666 -4098
rect 8853 -4174 15036 -4169
rect 8853 -4274 10700 -4174
rect 10764 -4274 15036 -4174
rect 8853 -4279 15036 -4274
rect 10674 -4408 10789 -4403
rect 10674 -4508 10700 -4408
rect 10764 -4508 10789 -4408
rect 10674 -4513 10789 -4508
rect 14926 -4579 15036 -4279
rect 6814 -4584 15036 -4579
rect 6814 -4684 6824 -4584
rect 6888 -4684 14576 -4584
rect 14640 -4684 15036 -4584
rect 6814 -4689 15036 -4684
<< via3 >>
rect 6813 1029 6877 2029
rect 8566 1029 8630 2029
rect 15543 443 15607 4467
rect 7690 -2132 7754 -1132
rect 6824 -4098 6888 -3998
rect 14593 -1665 14657 -1545
rect 14592 -2541 14656 -2421
rect 14576 -4098 14640 -3998
rect 10700 -4508 10764 -4408
<< mimcap >>
rect 11295 4415 15295 4455
rect 11295 495 11335 4415
rect 15255 495 15295 4415
rect 11295 455 15295 495
<< mimcapcontact >>
rect 11335 495 15255 4415
<< metal4 >>
rect 15527 4467 15623 4483
rect 11334 4415 15256 4416
rect 6812 2029 6878 2030
rect 6812 1029 6813 2029
rect 6877 1128 6878 2029
rect 8565 2029 8631 2030
rect 8565 1128 8566 2029
rect 6877 1029 8566 1128
rect 8630 1128 8631 2029
rect 8630 1029 9266 1128
rect 6812 1028 9266 1029
rect 7689 -1132 7755 -1131
rect 7689 -2132 7690 -1132
rect 7754 -1166 7755 -1132
rect 9166 -1166 9266 1028
rect 11334 495 11335 4415
rect 15255 495 15256 4415
rect 11334 494 15256 495
rect 7754 -1266 9266 -1166
rect 7754 -2132 7755 -1266
rect 7689 -2133 7755 -2132
rect 9166 -3997 9266 -1266
rect 14592 -1545 14658 494
rect 15527 443 15543 4467
rect 15607 443 15623 4467
rect 15527 427 15623 443
rect 14592 -1665 14593 -1545
rect 14657 -1665 14658 -1545
rect 14592 -1666 14658 -1665
rect 14591 -2421 14657 -2420
rect 14591 -2541 14592 -2421
rect 14656 -2541 14657 -2421
rect 14591 -3997 14657 -2541
rect 6823 -3998 15304 -3997
rect 6823 -4098 6824 -3998
rect 6888 -4098 14576 -3998
rect 14640 -4098 15304 -3998
rect 6823 -4099 15304 -4098
rect 15202 -4407 15304 -4099
rect 10699 -4408 15304 -4407
rect 10699 -4508 10700 -4408
rect 10764 -4508 15304 -4408
rect 10699 -4509 15304 -4508
<< labels >>
rlabel metal2 6403 4402 6403 4402 7 vcc
port 1 w
rlabel metal2 6498 -5017 6498 -5017 7 vss
port 2 w
rlabel metal4 15303 -4254 15303 -4254 3 vo
port 3 e
rlabel metal1 6297 687 6297 687 3 vd1
port 4 e
rlabel metal1 6297 372 6297 372 7 vd2
port 5 w
rlabel metal2 15099 -5082 15099 -5082 5 vb1
port 6 s
<< end >>
