VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DalinEM_diff_amp
  CLASS BLOCK ;
  FOREIGN tt_um_DalinEM_diff_amp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.524000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 144.000000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 144.000000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 15.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 74.780495 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 157.000 5.000 159.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.000 5.000 4.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 52.115 37.675 67.685 48.465 ;
      LAYER nwell ;
        RECT 75.155 48.375 78.315 48.395 ;
      LAYER pwell ;
        RECT 67.915 47.430 74.615 48.195 ;
        RECT 67.915 42.260 68.680 47.430 ;
        RECT 73.850 42.260 74.615 47.430 ;
      LAYER nwell ;
        RECT 75.155 42.475 78.320 48.375 ;
      LAYER pwell ;
        RECT 67.915 41.495 74.615 42.260 ;
        RECT 52.115 37.665 58.585 37.675 ;
        RECT 52.115 37.505 58.335 37.665 ;
        RECT 58.355 37.510 58.585 37.665 ;
        RECT 58.600 37.510 67.685 37.675 ;
        RECT 58.355 37.505 67.685 37.510 ;
        RECT 52.115 14.255 67.685 37.505 ;
        RECT 70.660 10.290 74.895 38.660 ;
      LAYER nwell ;
        RECT 75.160 38.320 78.320 42.475 ;
        RECT 75.120 32.645 78.310 36.605 ;
        RECT 75.120 26.195 78.310 30.155 ;
        RECT 108.880 26.560 148.930 33.935 ;
        RECT 75.120 19.745 78.310 23.705 ;
        RECT 75.200 10.360 78.375 17.225 ;
      LAYER pwell ;
        RECT 108.900 8.990 114.000 15.950 ;
        RECT 115.200 6.335 142.835 24.110 ;
        RECT 115.620 6.165 115.735 6.335 ;
        RECT 116.205 6.165 142.370 6.175 ;
      LAYER li1 ;
        RECT 77.810 48.585 79.980 48.590 ;
        RECT 51.740 48.055 53.545 48.490 ;
        RECT 77.810 48.205 80.160 48.585 ;
        RECT 68.045 48.060 74.485 48.065 ;
        RECT 67.615 48.055 74.485 48.060 ;
        RECT 51.740 47.595 74.485 48.055 ;
        RECT 51.740 15.480 53.545 47.595 ;
        RECT 66.610 46.890 74.485 47.595 ;
        RECT 54.175 46.695 58.215 46.865 ;
        RECT 61.580 46.695 65.620 46.865 ;
        RECT 66.610 46.795 69.220 46.890 ;
        RECT 53.835 45.635 54.005 46.635 ;
        RECT 58.385 45.635 58.555 46.635 ;
        RECT 61.240 45.635 61.410 46.635 ;
        RECT 65.790 45.635 65.960 46.635 ;
        RECT 54.175 45.405 58.215 45.575 ;
        RECT 61.580 45.405 65.620 45.575 ;
        RECT 53.835 44.345 54.005 45.345 ;
        RECT 58.385 44.345 58.555 45.345 ;
        RECT 61.240 44.345 61.410 45.345 ;
        RECT 65.790 44.345 65.960 45.345 ;
        RECT 54.175 44.115 58.215 44.285 ;
        RECT 61.580 44.115 65.620 44.285 ;
        RECT 53.835 43.055 54.005 44.055 ;
        RECT 58.385 43.055 58.555 44.055 ;
        RECT 61.240 43.055 61.410 44.055 ;
        RECT 65.790 43.055 65.960 44.055 ;
        RECT 54.175 42.825 58.215 42.995 ;
        RECT 61.580 42.825 65.620 42.995 ;
        RECT 66.575 42.800 69.220 46.795 ;
        RECT 69.530 43.110 73.000 46.580 ;
        RECT 73.310 42.800 74.485 46.890 ;
        RECT 53.835 41.765 54.005 42.765 ;
        RECT 58.385 41.765 58.555 42.765 ;
        RECT 61.240 41.765 61.410 42.765 ;
        RECT 65.790 41.765 65.960 42.765 ;
        RECT 54.175 41.535 58.215 41.705 ;
        RECT 61.580 41.535 65.620 41.705 ;
        RECT 66.575 41.625 74.485 42.800 ;
        RECT 75.350 47.945 80.160 48.205 ;
        RECT 53.835 40.475 54.005 41.475 ;
        RECT 58.385 40.475 58.555 41.475 ;
        RECT 61.240 40.475 61.410 41.475 ;
        RECT 65.790 40.475 65.960 41.475 ;
        RECT 54.175 40.245 58.215 40.415 ;
        RECT 61.580 40.245 65.620 40.415 ;
        RECT 53.835 39.185 54.005 40.185 ;
        RECT 58.385 39.185 58.555 40.185 ;
        RECT 61.240 39.185 61.410 40.185 ;
        RECT 65.790 39.185 65.960 40.185 ;
        RECT 54.175 38.955 58.215 39.125 ;
        RECT 61.580 38.955 65.620 39.125 ;
        RECT 53.835 37.895 54.005 38.895 ;
        RECT 58.385 37.895 58.555 38.895 ;
        RECT 61.240 37.895 61.410 38.895 ;
        RECT 65.790 37.895 65.960 38.895 ;
        RECT 66.575 38.510 68.075 41.625 ;
        RECT 75.350 38.745 75.590 47.945 ;
        RECT 76.200 47.285 76.740 47.455 ;
        RECT 77.810 47.390 80.160 47.945 ;
        RECT 75.815 45.225 75.985 47.225 ;
        RECT 76.955 45.225 77.125 47.225 ;
        RECT 77.815 47.160 80.160 47.390 ;
        RECT 76.200 44.995 76.740 45.165 ;
        RECT 75.815 42.935 75.985 44.935 ;
        RECT 76.955 42.935 77.125 44.935 ;
        RECT 76.200 42.705 76.740 42.875 ;
        RECT 77.810 42.220 80.160 47.160 ;
        RECT 76.200 41.660 77.240 41.830 ;
        RECT 75.815 40.600 75.985 41.600 ;
        RECT 77.455 40.600 77.625 41.600 ;
        RECT 76.200 40.370 77.240 40.540 ;
        RECT 75.815 39.310 75.985 40.310 ;
        RECT 77.455 39.310 77.625 40.310 ;
        RECT 76.200 39.080 77.240 39.250 ;
        RECT 77.825 38.905 80.160 42.220 ;
        RECT 77.495 38.745 80.160 38.905 ;
        RECT 66.575 38.505 70.445 38.510 ;
        RECT 66.575 37.890 74.850 38.505 ;
        RECT 75.350 38.500 80.160 38.745 ;
        RECT 54.175 37.665 58.215 37.835 ;
        RECT 61.580 37.665 65.620 37.835 ;
        RECT 53.835 36.605 54.005 37.605 ;
        RECT 58.385 36.605 58.555 37.605 ;
        RECT 61.240 36.605 61.410 37.605 ;
        RECT 65.790 36.605 65.960 37.605 ;
        RECT 54.175 36.375 58.215 36.545 ;
        RECT 61.580 36.375 65.620 36.545 ;
        RECT 53.835 35.315 54.005 36.315 ;
        RECT 58.385 35.315 58.555 36.315 ;
        RECT 61.240 35.315 61.410 36.315 ;
        RECT 65.790 35.315 65.960 36.315 ;
        RECT 54.175 35.085 58.215 35.255 ;
        RECT 61.580 35.085 65.620 35.255 ;
        RECT 53.835 34.025 54.005 35.025 ;
        RECT 58.385 34.025 58.555 35.025 ;
        RECT 61.240 34.025 61.410 35.025 ;
        RECT 65.790 34.025 65.960 35.025 ;
        RECT 54.175 33.795 58.215 33.965 ;
        RECT 61.580 33.795 65.620 33.965 ;
        RECT 53.835 32.735 54.005 33.735 ;
        RECT 58.385 32.735 58.555 33.735 ;
        RECT 61.240 32.735 61.410 33.735 ;
        RECT 65.790 32.735 65.960 33.735 ;
        RECT 54.175 32.505 58.215 32.675 ;
        RECT 61.580 32.505 65.620 32.675 ;
        RECT 53.835 31.445 54.005 32.445 ;
        RECT 58.385 31.445 58.555 32.445 ;
        RECT 61.240 31.445 61.410 32.445 ;
        RECT 65.790 31.445 65.960 32.445 ;
        RECT 54.175 31.215 58.215 31.385 ;
        RECT 61.580 31.215 65.620 31.385 ;
        RECT 53.835 30.155 54.005 31.155 ;
        RECT 58.385 30.155 58.555 31.155 ;
        RECT 61.240 30.155 61.410 31.155 ;
        RECT 65.790 30.155 65.960 31.155 ;
        RECT 54.175 29.925 58.215 30.095 ;
        RECT 61.580 29.925 65.620 30.095 ;
        RECT 53.835 28.865 54.005 29.865 ;
        RECT 58.385 28.865 58.555 29.865 ;
        RECT 61.240 28.865 61.410 29.865 ;
        RECT 65.790 28.865 65.960 29.865 ;
        RECT 54.175 28.635 58.215 28.805 ;
        RECT 61.580 28.635 65.620 28.805 ;
        RECT 53.835 27.575 54.005 28.575 ;
        RECT 58.385 27.575 58.555 28.575 ;
        RECT 61.240 27.575 61.410 28.575 ;
        RECT 65.790 27.575 65.960 28.575 ;
        RECT 54.175 27.345 58.215 27.515 ;
        RECT 61.580 27.345 65.620 27.515 ;
        RECT 53.835 26.285 54.005 27.285 ;
        RECT 58.385 26.285 58.555 27.285 ;
        RECT 61.240 26.285 61.410 27.285 ;
        RECT 65.790 26.285 65.960 27.285 ;
        RECT 54.175 26.055 58.215 26.225 ;
        RECT 61.580 26.055 65.620 26.225 ;
        RECT 53.835 24.995 54.005 25.995 ;
        RECT 58.385 24.995 58.555 25.995 ;
        RECT 61.240 24.995 61.410 25.995 ;
        RECT 65.790 24.995 65.960 25.995 ;
        RECT 54.175 24.765 58.215 24.935 ;
        RECT 61.580 24.765 65.620 24.935 ;
        RECT 53.835 23.705 54.005 24.705 ;
        RECT 58.385 23.705 58.555 24.705 ;
        RECT 61.240 23.705 61.410 24.705 ;
        RECT 65.790 23.705 65.960 24.705 ;
        RECT 54.175 23.475 58.215 23.645 ;
        RECT 61.580 23.475 65.620 23.645 ;
        RECT 53.835 22.415 54.005 23.415 ;
        RECT 58.385 22.415 58.555 23.415 ;
        RECT 61.240 22.415 61.410 23.415 ;
        RECT 65.790 22.415 65.960 23.415 ;
        RECT 54.175 22.185 58.215 22.355 ;
        RECT 61.580 22.185 65.620 22.355 ;
        RECT 53.835 21.125 54.005 22.125 ;
        RECT 58.385 21.125 58.555 22.125 ;
        RECT 61.240 21.125 61.410 22.125 ;
        RECT 65.790 21.125 65.960 22.125 ;
        RECT 54.175 20.895 58.215 21.065 ;
        RECT 61.580 20.895 65.620 21.065 ;
        RECT 53.835 19.835 54.005 20.835 ;
        RECT 58.385 19.835 58.555 20.835 ;
        RECT 61.240 19.835 61.410 20.835 ;
        RECT 65.790 19.835 65.960 20.835 ;
        RECT 54.175 19.605 58.215 19.775 ;
        RECT 61.580 19.605 65.620 19.775 ;
        RECT 53.835 18.545 54.005 19.545 ;
        RECT 58.385 18.545 58.555 19.545 ;
        RECT 61.240 18.545 61.410 19.545 ;
        RECT 65.790 18.545 65.960 19.545 ;
        RECT 54.175 18.315 58.215 18.485 ;
        RECT 61.580 18.315 65.620 18.485 ;
        RECT 53.835 17.255 54.005 18.255 ;
        RECT 58.385 17.255 58.555 18.255 ;
        RECT 61.240 17.255 61.410 18.255 ;
        RECT 65.790 17.255 65.960 18.255 ;
        RECT 54.175 17.025 58.215 17.195 ;
        RECT 61.580 17.025 65.620 17.195 ;
        RECT 53.835 15.965 54.005 16.965 ;
        RECT 58.385 15.965 58.555 16.965 ;
        RECT 61.240 15.965 61.410 16.965 ;
        RECT 65.790 15.965 65.960 16.965 ;
        RECT 54.175 15.735 58.215 15.905 ;
        RECT 61.580 15.735 65.620 15.905 ;
        RECT 66.575 15.480 71.680 37.890 ;
        RECT 72.260 37.265 73.300 37.435 ;
        RECT 71.920 36.205 72.090 37.205 ;
        RECT 73.470 36.205 73.640 37.205 ;
        RECT 72.260 35.975 73.300 36.145 ;
        RECT 71.920 34.915 72.090 35.915 ;
        RECT 73.470 34.915 73.640 35.915 ;
        RECT 72.260 34.685 73.300 34.855 ;
        RECT 71.920 33.625 72.090 34.625 ;
        RECT 73.470 33.625 73.640 34.625 ;
        RECT 72.260 33.395 73.300 33.565 ;
        RECT 71.920 32.335 72.090 33.335 ;
        RECT 73.470 32.335 73.640 33.335 ;
        RECT 72.260 32.105 73.300 32.275 ;
        RECT 71.920 31.045 72.090 32.045 ;
        RECT 73.470 31.045 73.640 32.045 ;
        RECT 72.260 30.815 73.300 30.985 ;
        RECT 71.920 29.755 72.090 30.755 ;
        RECT 73.470 29.755 73.640 30.755 ;
        RECT 72.260 29.525 73.300 29.695 ;
        RECT 71.920 28.465 72.090 29.465 ;
        RECT 73.470 28.465 73.640 29.465 ;
        RECT 72.260 28.235 73.300 28.405 ;
        RECT 71.920 27.175 72.090 28.175 ;
        RECT 73.470 27.175 73.640 28.175 ;
        RECT 72.260 26.945 73.300 27.115 ;
        RECT 71.920 25.885 72.090 26.885 ;
        RECT 73.470 25.885 73.640 26.885 ;
        RECT 72.260 25.655 73.300 25.825 ;
        RECT 71.920 24.595 72.090 25.595 ;
        RECT 73.470 24.595 73.640 25.595 ;
        RECT 72.260 24.365 73.300 24.535 ;
        RECT 71.920 23.305 72.090 24.305 ;
        RECT 73.470 23.305 73.640 24.305 ;
        RECT 72.260 23.075 73.300 23.245 ;
        RECT 71.920 22.015 72.090 23.015 ;
        RECT 73.470 22.015 73.640 23.015 ;
        RECT 72.260 21.785 73.300 21.955 ;
        RECT 71.920 20.725 72.090 21.725 ;
        RECT 73.470 20.725 73.640 21.725 ;
        RECT 72.260 20.495 73.300 20.665 ;
        RECT 71.920 19.435 72.090 20.435 ;
        RECT 73.470 19.435 73.640 20.435 ;
        RECT 72.260 19.205 73.300 19.375 ;
        RECT 71.920 18.145 72.090 19.145 ;
        RECT 73.470 18.145 73.640 19.145 ;
        RECT 72.260 17.915 73.300 18.085 ;
        RECT 71.920 16.855 72.090 17.855 ;
        RECT 73.470 16.855 73.640 17.855 ;
        RECT 72.260 16.625 73.300 16.795 ;
        RECT 71.920 15.565 72.090 16.565 ;
        RECT 73.470 15.565 73.640 16.565 ;
        RECT 51.740 14.900 71.680 15.480 ;
        RECT 72.260 15.335 73.300 15.505 ;
        RECT 70.400 11.010 71.680 14.900 ;
        RECT 71.920 14.275 72.090 15.275 ;
        RECT 73.470 14.275 73.640 15.275 ;
        RECT 72.260 14.045 73.300 14.215 ;
        RECT 71.920 12.985 72.090 13.985 ;
        RECT 73.470 12.985 73.640 13.985 ;
        RECT 72.260 12.755 73.300 12.925 ;
        RECT 71.920 11.695 72.090 12.695 ;
        RECT 73.470 11.695 73.640 12.695 ;
        RECT 72.260 11.465 73.300 11.635 ;
        RECT 74.155 11.010 74.850 37.890 ;
        RECT 77.495 38.285 80.160 38.500 ;
        RECT 77.495 36.540 80.150 38.285 ;
        RECT 75.200 36.530 80.150 36.540 ;
        RECT 75.190 36.150 80.150 36.530 ;
        RECT 75.190 33.090 75.530 36.150 ;
        RECT 77.495 36.135 80.150 36.150 ;
        RECT 76.195 35.685 77.235 35.855 ;
        RECT 75.810 33.625 75.980 35.625 ;
        RECT 77.450 33.625 77.620 35.625 ;
        RECT 76.195 33.395 77.235 33.565 ;
        RECT 77.860 33.090 80.150 36.135 ;
        RECT 75.190 32.700 80.150 33.090 ;
        RECT 75.190 32.695 75.530 32.700 ;
        RECT 75.220 30.125 75.600 30.145 ;
        RECT 76.110 30.125 80.150 32.700 ;
        RECT 75.220 29.700 80.150 30.125 ;
        RECT 75.220 26.595 75.600 29.700 ;
        RECT 76.195 29.235 77.235 29.405 ;
        RECT 75.810 27.175 75.980 29.175 ;
        RECT 77.450 27.175 77.620 29.175 ;
        RECT 76.195 26.945 77.235 27.115 ;
        RECT 77.860 26.595 80.150 29.700 ;
        RECT 75.220 26.195 80.150 26.595 ;
        RECT 108.350 32.865 149.230 34.555 ;
        RECT 108.350 27.020 109.620 32.865 ;
        RECT 110.825 32.420 128.825 32.590 ;
        RECT 129.115 32.420 147.115 32.590 ;
        RECT 110.595 30.365 110.765 32.205 ;
        RECT 128.885 30.365 129.055 32.205 ;
        RECT 147.175 30.365 147.345 32.205 ;
        RECT 110.825 29.980 128.825 30.150 ;
        RECT 129.115 29.980 147.115 30.150 ;
        RECT 110.595 27.925 110.765 29.765 ;
        RECT 128.885 27.925 129.055 29.765 ;
        RECT 147.175 27.925 147.345 29.765 ;
        RECT 110.825 27.540 128.825 27.710 ;
        RECT 129.115 27.540 147.115 27.710 ;
        RECT 148.180 27.020 149.225 32.865 ;
        RECT 108.350 26.355 149.225 27.020 ;
        RECT 76.050 23.665 80.150 26.195 ;
        RECT 75.175 23.210 80.150 23.665 ;
        RECT 75.175 20.225 75.590 23.210 ;
        RECT 76.195 22.785 77.235 22.955 ;
        RECT 77.855 22.730 80.150 23.210 ;
        RECT 75.810 20.725 75.980 22.725 ;
        RECT 77.450 20.725 77.620 22.725 ;
        RECT 76.195 20.495 77.235 20.665 ;
        RECT 77.860 20.230 80.150 22.730 ;
        RECT 77.855 20.225 80.150 20.230 ;
        RECT 75.175 19.745 80.150 20.225 ;
        RECT 76.050 17.205 80.150 19.745 ;
        RECT 75.230 17.195 80.150 17.205 ;
        RECT 70.400 10.395 74.850 11.010 ;
        RECT 75.220 16.780 80.150 17.195 ;
        RECT 75.220 10.865 75.615 16.780 ;
        RECT 76.195 16.335 77.235 16.505 ;
        RECT 75.810 14.275 75.980 16.275 ;
        RECT 77.450 14.275 77.620 16.275 ;
        RECT 76.195 14.045 77.235 14.215 ;
        RECT 76.195 13.430 77.235 13.600 ;
        RECT 75.810 11.370 75.980 13.370 ;
        RECT 77.450 11.370 77.620 13.370 ;
        RECT 76.195 11.140 77.235 11.310 ;
        RECT 77.860 10.865 80.150 16.780 ;
        RECT 108.355 23.480 144.100 24.180 ;
        RECT 108.355 15.775 115.735 23.480 ;
        RECT 116.875 23.015 128.875 23.185 ;
        RECT 129.165 23.015 141.165 23.185 ;
        RECT 116.645 16.805 116.815 22.845 ;
        RECT 128.935 16.805 129.105 22.845 ;
        RECT 141.225 16.805 141.395 22.845 ;
        RECT 116.875 16.465 128.875 16.635 ;
        RECT 129.165 16.465 141.165 16.635 ;
        RECT 75.220 10.350 80.150 10.865 ;
        RECT 75.220 10.345 77.940 10.350 ;
        RECT 79.360 10.315 80.150 10.350 ;
        RECT 108.350 15.590 115.735 15.775 ;
        RECT 108.350 9.360 109.405 15.590 ;
        RECT 109.930 15.030 112.970 15.200 ;
        RECT 109.590 9.970 109.760 14.970 ;
        RECT 113.140 9.970 113.310 14.970 ;
        RECT 109.930 9.360 112.970 9.910 ;
        RECT 113.610 9.360 115.735 15.590 ;
        RECT 116.870 13.640 128.870 13.810 ;
        RECT 129.160 13.640 141.160 13.810 ;
        RECT 108.350 8.210 115.735 9.360 ;
        RECT 108.340 6.810 115.735 8.210 ;
        RECT 116.640 7.430 116.810 13.470 ;
        RECT 128.930 7.430 129.100 13.470 ;
        RECT 141.220 7.430 141.390 13.470 ;
        RECT 116.870 7.090 128.870 7.260 ;
        RECT 129.160 7.090 141.160 7.260 ;
        RECT 142.350 6.810 144.100 23.480 ;
        RECT 108.340 5.260 144.100 6.810 ;
      LAYER met1 ;
        RECT 52.100 15.025 53.030 48.035 ;
        RECT 53.410 47.990 54.170 48.010 ;
        RECT 58.360 47.990 59.100 48.010 ;
        RECT 53.350 47.660 54.230 47.990 ;
        RECT 58.300 47.660 59.160 47.990 ;
        RECT 70.700 47.810 73.095 47.830 ;
        RECT 53.410 47.640 54.170 47.660 ;
        RECT 58.360 47.640 59.100 47.660 ;
        RECT 59.470 47.280 70.000 47.540 ;
        RECT 54.255 46.895 55.255 46.990 ;
        RECT 54.195 46.665 58.195 46.895 ;
        RECT 53.805 46.370 54.035 46.615 ;
        RECT 54.255 46.570 55.255 46.665 ;
        RECT 58.355 46.370 58.585 46.615 ;
        RECT 53.805 45.925 58.585 46.370 ;
        RECT 53.805 45.050 54.035 45.925 ;
        RECT 57.135 45.605 58.135 45.680 ;
        RECT 54.195 45.375 58.195 45.605 ;
        RECT 57.135 45.300 58.135 45.375 ;
        RECT 58.355 45.050 58.585 45.925 ;
        RECT 53.805 44.975 58.585 45.050 ;
        RECT 53.805 44.605 58.600 44.975 ;
        RECT 53.805 44.365 54.035 44.605 ;
        RECT 56.015 44.315 56.515 44.380 ;
        RECT 58.340 44.375 58.600 44.605 ;
        RECT 58.355 44.365 58.585 44.375 ;
        RECT 54.195 44.085 58.195 44.315 ;
        RECT 53.805 43.805 54.035 44.035 ;
        RECT 56.015 44.020 56.515 44.085 ;
        RECT 58.355 43.805 58.585 44.035 ;
        RECT 53.805 43.360 58.585 43.805 ;
        RECT 53.805 42.485 54.035 43.360 ;
        RECT 54.255 43.025 55.255 43.090 ;
        RECT 54.195 42.795 58.195 43.025 ;
        RECT 54.255 42.730 55.255 42.795 ;
        RECT 58.355 42.485 58.585 43.360 ;
        RECT 53.805 42.395 58.585 42.485 ;
        RECT 53.805 42.045 58.600 42.395 ;
        RECT 53.805 41.785 54.035 42.045 ;
        RECT 56.015 41.735 56.515 41.800 ;
        RECT 58.340 41.795 58.600 42.045 ;
        RECT 58.355 41.785 58.585 41.795 ;
        RECT 54.195 41.505 58.195 41.735 ;
        RECT 53.805 41.180 54.035 41.455 ;
        RECT 56.015 41.440 56.515 41.505 ;
        RECT 58.355 41.180 58.585 41.455 ;
        RECT 53.805 40.740 58.585 41.180 ;
        RECT 53.805 39.865 54.035 40.740 ;
        RECT 57.135 40.445 58.135 40.520 ;
        RECT 54.195 40.215 58.195 40.445 ;
        RECT 57.135 40.140 58.135 40.215 ;
        RECT 58.355 39.865 58.585 40.740 ;
        RECT 53.805 39.425 58.585 39.865 ;
        RECT 53.805 38.615 54.035 39.425 ;
        RECT 54.255 39.155 55.255 39.250 ;
        RECT 54.195 38.925 58.195 39.155 ;
        RECT 54.255 38.830 55.255 38.925 ;
        RECT 58.355 38.615 58.585 39.425 ;
        RECT 53.805 38.175 58.585 38.615 ;
        RECT 53.805 37.320 54.035 38.175 ;
        RECT 57.135 37.865 58.135 37.940 ;
        RECT 54.195 37.635 58.195 37.865 ;
        RECT 57.135 37.560 58.135 37.635 ;
        RECT 58.355 37.430 58.585 38.175 ;
        RECT 58.290 37.320 58.650 37.430 ;
        RECT 53.805 37.205 58.650 37.320 ;
        RECT 53.805 36.880 58.600 37.205 ;
        RECT 53.805 36.625 54.035 36.880 ;
        RECT 56.015 36.575 56.515 36.640 ;
        RECT 58.340 36.635 58.600 36.880 ;
        RECT 58.355 36.625 58.585 36.635 ;
        RECT 54.195 36.345 58.195 36.575 ;
        RECT 53.805 36.055 54.035 36.295 ;
        RECT 56.015 36.280 56.515 36.345 ;
        RECT 58.355 36.055 58.585 36.295 ;
        RECT 53.805 35.590 58.585 36.055 ;
        RECT 53.805 34.745 54.035 35.590 ;
        RECT 54.255 35.285 55.255 35.350 ;
        RECT 54.195 35.055 58.195 35.285 ;
        RECT 54.255 34.990 55.255 35.055 ;
        RECT 58.355 34.745 58.585 35.590 ;
        RECT 53.805 34.655 58.585 34.745 ;
        RECT 53.805 34.305 58.600 34.655 ;
        RECT 53.805 34.045 54.035 34.305 ;
        RECT 56.015 33.995 56.515 34.060 ;
        RECT 58.340 34.055 58.600 34.305 ;
        RECT 58.355 34.045 58.585 34.055 ;
        RECT 54.195 33.765 58.195 33.995 ;
        RECT 53.805 33.420 54.035 33.715 ;
        RECT 56.015 33.700 56.515 33.765 ;
        RECT 58.355 33.420 58.585 33.715 ;
        RECT 53.805 32.980 58.585 33.420 ;
        RECT 53.805 32.140 54.035 32.980 ;
        RECT 57.135 32.705 58.135 32.780 ;
        RECT 54.195 32.475 58.195 32.705 ;
        RECT 57.135 32.400 58.135 32.475 ;
        RECT 58.355 32.140 58.585 32.980 ;
        RECT 53.805 31.700 58.585 32.140 ;
        RECT 53.805 30.855 54.035 31.700 ;
        RECT 54.255 31.415 55.255 31.510 ;
        RECT 54.195 31.185 58.195 31.415 ;
        RECT 54.255 31.090 55.255 31.185 ;
        RECT 58.355 30.855 58.585 31.700 ;
        RECT 53.805 30.415 58.585 30.855 ;
        RECT 53.805 29.560 54.035 30.415 ;
        RECT 57.135 30.125 58.135 30.200 ;
        RECT 54.195 29.895 58.195 30.125 ;
        RECT 57.135 29.820 58.135 29.895 ;
        RECT 58.355 29.645 58.585 30.415 ;
        RECT 58.340 29.560 58.600 29.645 ;
        RECT 53.805 29.120 58.600 29.560 ;
        RECT 53.805 28.885 54.035 29.120 ;
        RECT 56.015 28.835 56.515 28.900 ;
        RECT 58.340 28.895 58.600 29.120 ;
        RECT 58.355 28.885 58.585 28.895 ;
        RECT 54.195 28.605 58.195 28.835 ;
        RECT 53.805 28.300 54.035 28.555 ;
        RECT 56.015 28.540 56.515 28.605 ;
        RECT 58.355 28.300 58.585 28.555 ;
        RECT 53.805 27.860 58.585 28.300 ;
        RECT 53.805 27.015 54.035 27.860 ;
        RECT 54.255 27.545 55.255 27.615 ;
        RECT 54.195 27.315 58.195 27.545 ;
        RECT 54.255 27.255 55.255 27.315 ;
        RECT 58.355 27.015 58.585 27.860 ;
        RECT 53.805 26.915 58.585 27.015 ;
        RECT 53.805 26.575 58.600 26.915 ;
        RECT 53.805 26.305 54.035 26.575 ;
        RECT 56.015 26.255 56.515 26.320 ;
        RECT 58.340 26.315 58.600 26.575 ;
        RECT 58.355 26.305 58.585 26.315 ;
        RECT 54.195 26.025 58.195 26.255 ;
        RECT 53.805 25.680 54.035 25.975 ;
        RECT 56.015 25.960 56.515 26.025 ;
        RECT 58.355 25.680 58.585 25.975 ;
        RECT 53.805 25.240 58.585 25.680 ;
        RECT 53.805 24.460 54.035 25.240 ;
        RECT 57.135 24.965 58.135 25.040 ;
        RECT 54.195 24.735 58.195 24.965 ;
        RECT 57.135 24.660 58.135 24.735 ;
        RECT 58.355 24.460 58.585 25.240 ;
        RECT 53.805 24.020 58.585 24.460 ;
        RECT 53.805 23.135 54.035 24.020 ;
        RECT 54.255 23.675 55.255 23.770 ;
        RECT 54.195 23.445 58.195 23.675 ;
        RECT 54.255 23.350 55.255 23.445 ;
        RECT 58.355 23.135 58.585 24.020 ;
        RECT 53.805 22.695 58.585 23.135 ;
        RECT 53.805 21.880 54.035 22.695 ;
        RECT 57.135 22.385 58.135 22.460 ;
        RECT 54.195 22.155 58.195 22.385 ;
        RECT 57.135 22.080 58.135 22.155 ;
        RECT 58.355 21.880 58.585 22.695 ;
        RECT 53.805 21.860 58.585 21.880 ;
        RECT 53.805 21.440 58.600 21.860 ;
        RECT 53.805 21.145 54.035 21.440 ;
        RECT 56.015 21.095 56.515 21.160 ;
        RECT 58.340 21.155 58.600 21.440 ;
        RECT 58.355 21.145 58.585 21.155 ;
        RECT 54.195 20.865 58.195 21.095 ;
        RECT 53.805 20.550 54.035 20.815 ;
        RECT 56.015 20.800 56.515 20.865 ;
        RECT 58.355 20.550 58.585 20.815 ;
        RECT 53.805 20.110 58.585 20.550 ;
        RECT 53.805 19.265 54.035 20.110 ;
        RECT 54.255 19.805 55.255 19.870 ;
        RECT 54.195 19.575 58.195 19.805 ;
        RECT 54.255 19.510 55.255 19.575 ;
        RECT 58.355 19.265 58.585 20.110 ;
        RECT 53.805 19.175 58.585 19.265 ;
        RECT 53.805 18.825 58.600 19.175 ;
        RECT 53.805 18.565 54.035 18.825 ;
        RECT 56.015 18.515 56.515 18.580 ;
        RECT 58.340 18.575 58.600 18.825 ;
        RECT 58.355 18.565 58.585 18.575 ;
        RECT 54.195 18.285 58.195 18.515 ;
        RECT 53.805 17.895 54.035 18.235 ;
        RECT 56.015 18.220 56.515 18.285 ;
        RECT 58.355 17.895 58.585 18.235 ;
        RECT 53.805 17.455 58.585 17.895 ;
        RECT 53.805 16.680 54.035 17.455 ;
        RECT 57.135 17.225 58.135 17.300 ;
        RECT 54.195 16.995 58.195 17.225 ;
        RECT 57.135 16.920 58.135 16.995 ;
        RECT 58.355 16.680 58.585 17.455 ;
        RECT 53.805 16.595 58.585 16.680 ;
        RECT 53.805 16.240 58.600 16.595 ;
        RECT 53.805 15.985 54.035 16.240 ;
        RECT 54.255 15.935 55.255 16.030 ;
        RECT 58.340 15.995 58.600 16.240 ;
        RECT 58.355 15.985 58.585 15.995 ;
        RECT 54.195 15.705 58.195 15.935 ;
        RECT 59.470 15.755 59.730 47.280 ;
        RECT 64.540 46.895 65.540 46.960 ;
        RECT 61.600 46.665 65.600 46.895 ;
        RECT 60.195 15.755 60.455 46.585 ;
        RECT 61.210 46.330 61.440 46.615 ;
        RECT 64.540 46.600 65.540 46.665 ;
        RECT 65.760 46.330 65.990 46.615 ;
        RECT 61.210 46.265 65.990 46.330 ;
        RECT 61.195 45.890 65.990 46.265 ;
        RECT 61.195 45.665 61.455 45.890 ;
        RECT 61.210 45.655 61.440 45.665 ;
        RECT 63.165 45.605 63.665 45.670 ;
        RECT 65.760 45.655 65.990 45.890 ;
        RECT 61.600 45.375 65.600 45.605 ;
        RECT 61.210 45.070 61.440 45.325 ;
        RECT 63.165 45.310 63.665 45.375 ;
        RECT 65.760 45.070 65.990 45.325 ;
        RECT 61.210 44.630 65.990 45.070 ;
        RECT 61.210 43.825 61.440 44.630 ;
        RECT 64.535 44.315 65.535 44.390 ;
        RECT 61.600 44.085 65.600 44.315 ;
        RECT 64.535 44.010 65.535 44.085 ;
        RECT 65.760 43.825 65.990 44.630 ;
        RECT 61.210 43.385 65.990 43.825 ;
        RECT 61.210 42.475 61.440 43.385 ;
        RECT 61.660 43.025 62.660 43.120 ;
        RECT 61.600 42.795 65.600 43.025 ;
        RECT 61.660 42.700 62.660 42.795 ;
        RECT 65.760 42.475 65.990 43.385 ;
        RECT 61.210 42.035 65.990 42.475 ;
        RECT 61.210 41.605 61.440 42.035 ;
        RECT 64.540 41.735 65.540 41.810 ;
        RECT 61.195 41.230 61.455 41.605 ;
        RECT 61.600 41.505 65.600 41.735 ;
        RECT 64.540 41.430 65.540 41.505 ;
        RECT 65.760 41.230 65.990 42.035 ;
        RECT 61.195 40.790 65.990 41.230 ;
        RECT 61.195 40.505 61.455 40.790 ;
        RECT 61.210 40.495 61.440 40.505 ;
        RECT 63.165 40.445 63.665 40.510 ;
        RECT 65.760 40.495 65.990 40.790 ;
        RECT 61.600 40.215 65.600 40.445 ;
        RECT 61.210 39.915 61.440 40.165 ;
        RECT 63.165 40.150 63.665 40.215 ;
        RECT 65.760 39.915 65.990 40.165 ;
        RECT 61.210 39.475 65.990 39.915 ;
        RECT 61.210 38.645 61.440 39.475 ;
        RECT 64.540 39.155 65.540 39.220 ;
        RECT 61.600 38.925 65.600 39.155 ;
        RECT 64.540 38.860 65.540 38.925 ;
        RECT 65.760 38.645 65.990 39.475 ;
        RECT 61.210 38.525 65.990 38.645 ;
        RECT 61.195 38.205 65.990 38.525 ;
        RECT 61.195 37.925 61.455 38.205 ;
        RECT 61.210 37.915 61.440 37.925 ;
        RECT 63.165 37.865 63.665 37.930 ;
        RECT 65.760 37.915 65.990 38.205 ;
        RECT 61.600 37.635 65.600 37.865 ;
        RECT 61.210 37.310 61.440 37.585 ;
        RECT 63.165 37.570 63.665 37.635 ;
        RECT 65.760 37.310 65.990 37.585 ;
        RECT 61.210 36.870 65.990 37.310 ;
        RECT 61.210 36.045 61.440 36.870 ;
        RECT 64.540 36.575 65.540 36.650 ;
        RECT 61.600 36.345 65.600 36.575 ;
        RECT 64.540 36.270 65.540 36.345 ;
        RECT 65.760 36.045 65.990 36.870 ;
        RECT 61.210 35.605 65.990 36.045 ;
        RECT 61.210 34.785 61.440 35.605 ;
        RECT 61.660 35.285 62.660 35.380 ;
        RECT 61.600 35.055 65.600 35.285 ;
        RECT 61.660 34.960 62.660 35.055 ;
        RECT 65.760 34.785 65.990 35.605 ;
        RECT 61.210 34.345 65.990 34.785 ;
        RECT 61.210 33.785 61.440 34.345 ;
        RECT 64.540 33.995 65.540 34.070 ;
        RECT 61.195 33.430 61.455 33.785 ;
        RECT 61.600 33.765 65.600 33.995 ;
        RECT 64.540 33.690 65.540 33.765 ;
        RECT 65.760 33.430 65.990 34.345 ;
        RECT 61.195 32.990 65.990 33.430 ;
        RECT 61.195 32.765 61.455 32.990 ;
        RECT 61.210 32.755 61.440 32.765 ;
        RECT 63.165 32.705 63.665 32.770 ;
        RECT 65.760 32.755 65.990 32.990 ;
        RECT 61.600 32.475 65.600 32.705 ;
        RECT 61.210 32.200 61.440 32.425 ;
        RECT 63.165 32.410 63.665 32.475 ;
        RECT 65.760 32.200 65.990 32.425 ;
        RECT 61.210 31.795 65.990 32.200 ;
        RECT 61.210 30.900 61.440 31.795 ;
        RECT 64.540 31.415 65.540 31.480 ;
        RECT 61.600 31.185 65.600 31.415 ;
        RECT 64.540 31.120 65.540 31.185 ;
        RECT 65.760 30.900 65.990 31.795 ;
        RECT 61.210 30.785 65.990 30.900 ;
        RECT 61.195 30.495 65.990 30.785 ;
        RECT 61.195 30.185 61.455 30.495 ;
        RECT 61.210 30.175 61.440 30.185 ;
        RECT 63.160 30.125 63.660 30.190 ;
        RECT 65.760 30.175 65.990 30.495 ;
        RECT 61.600 29.895 65.600 30.125 ;
        RECT 61.210 29.590 61.440 29.845 ;
        RECT 63.160 29.830 63.660 29.895 ;
        RECT 65.760 29.590 65.990 29.845 ;
        RECT 61.210 29.150 65.990 29.590 ;
        RECT 61.210 28.310 61.440 29.150 ;
        RECT 64.540 28.835 65.540 28.910 ;
        RECT 61.600 28.605 65.600 28.835 ;
        RECT 64.540 28.530 65.540 28.605 ;
        RECT 65.760 28.310 65.990 29.150 ;
        RECT 61.210 27.870 65.990 28.310 ;
        RECT 61.210 27.005 61.440 27.870 ;
        RECT 61.660 27.545 62.660 27.640 ;
        RECT 61.600 27.315 65.600 27.545 ;
        RECT 61.660 27.220 62.660 27.315 ;
        RECT 65.760 27.005 65.990 27.870 ;
        RECT 61.210 26.565 65.990 27.005 ;
        RECT 61.210 26.045 61.440 26.565 ;
        RECT 64.540 26.255 65.540 26.330 ;
        RECT 61.195 25.730 61.455 26.045 ;
        RECT 61.600 26.025 65.600 26.255 ;
        RECT 64.540 25.950 65.540 26.025 ;
        RECT 65.760 25.730 65.990 26.565 ;
        RECT 61.195 25.290 65.990 25.730 ;
        RECT 61.195 25.025 61.455 25.290 ;
        RECT 61.210 25.015 61.440 25.025 ;
        RECT 63.165 24.965 63.665 25.030 ;
        RECT 65.760 25.015 65.990 25.290 ;
        RECT 61.600 24.735 65.600 24.965 ;
        RECT 61.210 24.455 61.440 24.685 ;
        RECT 63.165 24.670 63.665 24.735 ;
        RECT 65.760 24.455 65.990 24.685 ;
        RECT 61.210 23.925 65.990 24.455 ;
        RECT 61.210 23.180 61.440 23.925 ;
        RECT 64.540 23.675 65.540 23.740 ;
        RECT 61.600 23.445 65.600 23.675 ;
        RECT 64.540 23.380 65.540 23.445 ;
        RECT 65.760 23.180 65.990 23.925 ;
        RECT 61.210 23.045 65.990 23.180 ;
        RECT 61.195 22.650 65.990 23.045 ;
        RECT 61.195 22.445 61.455 22.650 ;
        RECT 61.210 22.435 61.440 22.445 ;
        RECT 63.165 22.385 63.665 22.450 ;
        RECT 65.760 22.435 65.990 22.650 ;
        RECT 61.600 22.155 65.600 22.385 ;
        RECT 61.210 21.830 61.440 22.105 ;
        RECT 63.165 22.090 63.665 22.155 ;
        RECT 65.760 21.830 65.990 22.105 ;
        RECT 61.210 21.390 65.990 21.830 ;
        RECT 61.210 20.550 61.440 21.390 ;
        RECT 64.540 21.095 65.540 21.170 ;
        RECT 61.600 20.865 65.600 21.095 ;
        RECT 64.540 20.790 65.540 20.865 ;
        RECT 65.760 20.550 65.990 21.390 ;
        RECT 61.210 20.110 65.990 20.550 ;
        RECT 61.210 19.255 61.440 20.110 ;
        RECT 61.660 19.805 62.660 19.900 ;
        RECT 61.600 19.575 65.600 19.805 ;
        RECT 61.660 19.480 62.660 19.575 ;
        RECT 65.760 19.255 65.990 20.110 ;
        RECT 61.210 18.815 65.990 19.255 ;
        RECT 61.210 18.305 61.440 18.815 ;
        RECT 64.540 18.515 65.540 18.590 ;
        RECT 61.195 17.955 61.455 18.305 ;
        RECT 61.600 18.285 65.600 18.515 ;
        RECT 64.540 18.210 65.540 18.285 ;
        RECT 65.760 17.955 65.990 18.815 ;
        RECT 61.195 17.515 65.990 17.955 ;
        RECT 61.195 17.285 61.455 17.515 ;
        RECT 61.210 17.275 61.440 17.285 ;
        RECT 63.165 17.225 63.665 17.290 ;
        RECT 65.760 17.275 65.990 17.515 ;
        RECT 61.600 16.995 65.600 17.225 ;
        RECT 61.210 16.690 61.440 16.945 ;
        RECT 63.165 16.930 63.665 16.995 ;
        RECT 65.760 16.690 65.990 16.945 ;
        RECT 61.210 16.595 65.990 16.690 ;
        RECT 61.195 16.250 65.990 16.595 ;
        RECT 61.195 15.995 61.455 16.250 ;
        RECT 61.210 15.985 61.440 15.995 ;
        RECT 64.540 15.935 65.540 16.000 ;
        RECT 65.760 15.985 65.990 16.250 ;
        RECT 61.600 15.705 65.600 15.935 ;
        RECT 54.255 15.610 55.255 15.705 ;
        RECT 64.540 15.640 65.540 15.705 ;
        RECT 66.805 15.245 67.425 47.075 ;
        RECT 67.610 44.355 68.150 47.110 ;
        RECT 69.740 46.370 70.000 47.280 ;
        RECT 70.640 47.150 73.155 47.810 ;
        RECT 70.700 47.130 73.095 47.150 ;
        RECT 69.740 43.320 72.790 46.370 ;
        RECT 73.555 43.110 74.355 47.355 ;
        RECT 75.785 47.255 76.720 47.485 ;
        RECT 75.785 47.160 76.015 47.255 ;
        RECT 75.680 46.910 76.015 47.160 ;
        RECT 76.925 46.910 77.155 47.205 ;
        RECT 75.680 45.500 77.155 46.910 ;
        RECT 75.680 45.265 76.015 45.500 ;
        RECT 75.785 44.890 76.015 45.265 ;
        RECT 76.280 45.195 76.660 45.260 ;
        RECT 76.925 45.245 77.155 45.500 ;
        RECT 76.220 44.965 76.720 45.195 ;
        RECT 76.280 44.900 76.660 44.965 ;
        RECT 75.680 44.675 76.015 44.890 ;
        RECT 76.925 44.675 77.155 44.915 ;
        RECT 75.680 43.265 77.155 44.675 ;
        RECT 77.925 43.435 78.645 48.400 ;
        RECT 75.680 42.995 76.015 43.265 ;
        RECT 75.785 42.905 76.015 42.995 ;
        RECT 76.925 42.955 77.155 43.265 ;
        RECT 75.785 42.675 76.720 42.905 ;
        RECT 68.535 42.575 73.750 42.595 ;
        RECT 68.475 41.975 73.810 42.575 ;
        RECT 68.535 41.955 73.750 41.975 ;
        RECT 75.785 41.365 76.015 42.675 ;
        RECT 76.280 41.860 76.980 41.955 ;
        RECT 76.220 41.630 77.220 41.860 ;
        RECT 76.280 41.535 76.980 41.630 ;
        RECT 77.425 41.365 77.655 41.580 ;
        RECT 75.785 40.775 77.655 41.365 ;
        RECT 75.785 40.105 76.015 40.775 ;
        RECT 76.460 40.570 77.160 40.635 ;
        RECT 77.425 40.620 77.655 40.775 ;
        RECT 76.220 40.340 77.220 40.570 ;
        RECT 76.460 40.275 77.160 40.340 ;
        RECT 77.425 40.105 77.655 40.290 ;
        RECT 75.785 39.695 77.655 40.105 ;
        RECT 75.780 39.515 77.655 39.695 ;
        RECT 70.510 10.945 71.525 38.100 ;
        RECT 72.340 37.465 72.640 37.530 ;
        RECT 72.280 37.235 73.280 37.465 ;
        RECT 71.890 36.880 72.120 37.185 ;
        RECT 72.340 37.170 72.640 37.235 ;
        RECT 73.440 36.880 73.670 37.185 ;
        RECT 71.890 36.545 73.670 36.880 ;
        RECT 71.890 35.590 72.120 36.545 ;
        RECT 72.340 36.175 72.640 36.240 ;
        RECT 72.280 35.945 73.280 36.175 ;
        RECT 72.340 35.880 72.640 35.945 ;
        RECT 73.440 35.590 73.670 36.545 ;
        RECT 71.890 35.255 73.670 35.590 ;
        RECT 71.890 34.885 72.120 35.255 ;
        RECT 73.440 34.950 73.670 35.255 ;
        RECT 72.920 34.885 73.670 34.950 ;
        RECT 71.890 34.655 73.670 34.885 ;
        RECT 71.890 34.280 72.120 34.655 ;
        RECT 72.920 34.590 73.670 34.655 ;
        RECT 73.440 34.280 73.670 34.590 ;
        RECT 71.890 33.945 73.670 34.280 ;
        RECT 71.890 32.995 72.120 33.945 ;
        RECT 72.340 33.595 72.640 33.660 ;
        RECT 72.280 33.365 73.280 33.595 ;
        RECT 72.340 33.300 72.640 33.365 ;
        RECT 73.440 32.995 73.670 33.945 ;
        RECT 71.890 32.660 73.670 32.995 ;
        RECT 71.890 32.305 72.120 32.660 ;
        RECT 73.440 32.370 73.670 32.660 ;
        RECT 72.920 32.305 73.670 32.370 ;
        RECT 71.890 32.075 73.670 32.305 ;
        RECT 71.890 31.695 72.120 32.075 ;
        RECT 72.920 32.010 73.670 32.075 ;
        RECT 73.440 31.695 73.670 32.010 ;
        RECT 71.890 31.360 73.670 31.695 ;
        RECT 71.890 31.065 72.120 31.360 ;
        RECT 72.340 31.015 72.640 31.080 ;
        RECT 73.440 31.065 73.670 31.360 ;
        RECT 75.780 36.455 76.015 39.515 ;
        RECT 76.280 39.280 76.980 39.375 ;
        RECT 77.425 39.330 77.655 39.515 ;
        RECT 76.220 39.050 77.220 39.280 ;
        RECT 76.280 38.955 76.980 39.050 ;
        RECT 77.915 38.385 78.650 43.435 ;
        RECT 78.980 38.380 79.780 48.395 ;
        RECT 75.780 35.355 76.010 36.455 ;
        RECT 76.540 35.885 77.155 35.950 ;
        RECT 76.215 35.655 77.215 35.885 ;
        RECT 76.540 35.590 77.155 35.655 ;
        RECT 77.420 35.355 77.650 35.605 ;
        RECT 75.780 33.960 77.650 35.355 ;
        RECT 72.280 30.785 73.280 31.015 ;
        RECT 71.890 30.435 72.120 30.735 ;
        RECT 72.340 30.720 72.640 30.785 ;
        RECT 73.440 30.435 73.670 30.735 ;
        RECT 71.890 30.100 73.670 30.435 ;
        RECT 71.890 29.165 72.120 30.100 ;
        RECT 72.340 29.725 72.640 29.790 ;
        RECT 72.280 29.495 73.280 29.725 ;
        RECT 72.340 29.430 72.640 29.495 ;
        RECT 73.440 29.165 73.670 30.100 ;
        RECT 71.890 28.830 73.670 29.165 ;
        RECT 71.890 28.435 72.120 28.830 ;
        RECT 73.440 28.500 73.670 28.830 ;
        RECT 72.920 28.435 73.670 28.500 ;
        RECT 71.890 28.205 73.670 28.435 ;
        RECT 71.890 27.860 72.120 28.205 ;
        RECT 72.920 28.140 73.670 28.205 ;
        RECT 73.440 27.860 73.670 28.140 ;
        RECT 71.890 27.525 73.670 27.860 ;
        RECT 71.890 26.595 72.120 27.525 ;
        RECT 72.340 27.145 72.640 27.210 ;
        RECT 72.280 26.915 73.280 27.145 ;
        RECT 72.340 26.850 72.640 26.915 ;
        RECT 73.440 26.595 73.670 27.525 ;
        RECT 71.890 26.260 73.670 26.595 ;
        RECT 71.890 25.855 72.120 26.260 ;
        RECT 73.440 25.920 73.670 26.260 ;
        RECT 72.920 25.855 73.670 25.920 ;
        RECT 71.890 25.625 73.670 25.855 ;
        RECT 71.890 25.285 72.120 25.625 ;
        RECT 72.920 25.560 73.670 25.625 ;
        RECT 73.440 25.285 73.670 25.560 ;
        RECT 71.890 24.950 73.670 25.285 ;
        RECT 71.890 24.615 72.120 24.950 ;
        RECT 72.340 24.565 72.640 24.630 ;
        RECT 73.440 24.615 73.670 24.950 ;
        RECT 75.780 28.865 76.010 33.960 ;
        RECT 76.275 33.595 76.840 33.660 ;
        RECT 77.420 33.645 77.650 33.960 ;
        RECT 76.215 33.365 77.215 33.595 ;
        RECT 76.275 33.300 76.840 33.365 ;
        RECT 76.540 29.435 77.155 29.500 ;
        RECT 76.215 29.205 77.215 29.435 ;
        RECT 76.540 29.140 77.155 29.205 ;
        RECT 77.420 28.865 77.650 29.155 ;
        RECT 75.780 27.470 77.650 28.865 ;
        RECT 72.280 24.335 73.280 24.565 ;
        RECT 71.890 23.995 72.120 24.285 ;
        RECT 72.340 24.270 72.640 24.335 ;
        RECT 73.440 23.995 73.670 24.285 ;
        RECT 71.890 23.660 73.670 23.995 ;
        RECT 71.890 22.710 72.120 23.660 ;
        RECT 72.340 23.275 72.640 23.340 ;
        RECT 72.280 23.045 73.280 23.275 ;
        RECT 72.340 22.980 72.640 23.045 ;
        RECT 73.440 22.710 73.670 23.660 ;
        RECT 71.890 22.375 73.670 22.710 ;
        RECT 71.890 21.985 72.120 22.375 ;
        RECT 73.440 22.050 73.670 22.375 ;
        RECT 72.920 21.985 73.670 22.050 ;
        RECT 71.890 21.755 73.670 21.985 ;
        RECT 71.890 21.405 72.120 21.755 ;
        RECT 72.920 21.690 73.670 21.755 ;
        RECT 73.440 21.405 73.670 21.690 ;
        RECT 71.890 21.070 73.670 21.405 ;
        RECT 71.890 20.110 72.120 21.070 ;
        RECT 72.340 20.695 72.640 20.760 ;
        RECT 72.280 20.465 73.280 20.695 ;
        RECT 72.340 20.400 72.640 20.465 ;
        RECT 73.440 20.110 73.670 21.070 ;
        RECT 71.890 19.775 73.670 20.110 ;
        RECT 71.890 19.405 72.120 19.775 ;
        RECT 73.440 19.470 73.670 19.775 ;
        RECT 72.920 19.405 73.670 19.470 ;
        RECT 71.890 19.175 73.670 19.405 ;
        RECT 71.890 18.860 72.120 19.175 ;
        RECT 72.920 19.110 73.670 19.175 ;
        RECT 73.440 18.860 73.670 19.110 ;
        RECT 71.890 18.525 73.670 18.860 ;
        RECT 71.890 18.165 72.120 18.525 ;
        RECT 72.340 18.115 72.640 18.180 ;
        RECT 73.440 18.165 73.670 18.525 ;
        RECT 75.780 22.460 76.010 27.470 ;
        RECT 76.275 27.145 76.840 27.210 ;
        RECT 77.420 27.195 77.650 27.470 ;
        RECT 76.215 26.915 77.215 27.145 ;
        RECT 76.275 26.850 76.840 26.915 ;
        RECT 76.540 22.985 77.155 23.050 ;
        RECT 76.215 22.755 77.215 22.985 ;
        RECT 76.540 22.690 77.155 22.755 ;
        RECT 77.420 22.460 77.650 22.705 ;
        RECT 75.780 21.065 77.650 22.460 ;
        RECT 72.280 17.885 73.280 18.115 ;
        RECT 71.890 17.560 72.120 17.835 ;
        RECT 72.340 17.820 72.640 17.885 ;
        RECT 73.440 17.560 73.670 17.835 ;
        RECT 71.890 17.225 73.670 17.560 ;
        RECT 71.890 16.250 72.120 17.225 ;
        RECT 72.340 16.825 72.640 16.890 ;
        RECT 72.280 16.595 73.280 16.825 ;
        RECT 72.340 16.530 72.640 16.595 ;
        RECT 73.440 16.250 73.670 17.225 ;
        RECT 71.890 15.915 73.670 16.250 ;
        RECT 71.890 15.535 72.120 15.915 ;
        RECT 73.440 15.600 73.670 15.915 ;
        RECT 72.920 15.535 73.670 15.600 ;
        RECT 71.890 15.305 73.670 15.535 ;
        RECT 71.890 14.950 72.120 15.305 ;
        RECT 72.920 15.240 73.670 15.305 ;
        RECT 73.440 14.950 73.670 15.240 ;
        RECT 71.890 14.615 73.670 14.950 ;
        RECT 71.890 13.655 72.120 14.615 ;
        RECT 72.340 14.245 72.640 14.310 ;
        RECT 72.280 14.015 73.280 14.245 ;
        RECT 72.340 13.950 72.640 14.015 ;
        RECT 73.440 13.655 73.670 14.615 ;
        RECT 71.890 13.320 73.670 13.655 ;
        RECT 71.890 12.955 72.120 13.320 ;
        RECT 73.440 13.020 73.670 13.320 ;
        RECT 72.920 12.955 73.670 13.020 ;
        RECT 71.890 12.725 73.670 12.955 ;
        RECT 71.890 12.320 72.120 12.725 ;
        RECT 72.920 12.660 73.670 12.725 ;
        RECT 73.440 12.320 73.670 12.660 ;
        RECT 71.890 11.985 73.670 12.320 ;
        RECT 71.890 11.715 72.120 11.985 ;
        RECT 72.340 11.665 72.640 11.730 ;
        RECT 72.920 11.665 73.220 11.730 ;
        RECT 73.440 11.715 73.670 11.985 ;
        RECT 75.780 15.910 76.010 21.065 ;
        RECT 76.275 20.695 76.840 20.760 ;
        RECT 77.420 20.745 77.650 21.065 ;
        RECT 76.215 20.465 77.215 20.695 ;
        RECT 76.275 20.400 76.840 20.465 ;
        RECT 78.480 17.490 79.235 35.950 ;
        RECT 109.210 33.900 148.320 34.405 ;
        RECT 109.860 32.390 147.095 32.620 ;
        RECT 109.860 30.380 110.860 32.390 ;
        RECT 109.860 25.225 110.290 30.380 ;
        RECT 111.745 30.180 127.940 32.390 ;
        RECT 128.855 32.125 129.085 32.185 ;
        RECT 128.785 30.445 129.155 32.125 ;
        RECT 128.855 30.385 129.085 30.445 ;
        RECT 130.055 30.180 146.250 32.390 ;
        RECT 147.075 30.390 148.085 32.190 ;
        RECT 147.145 30.385 147.375 30.390 ;
        RECT 110.845 29.950 128.805 30.180 ;
        RECT 129.135 29.950 147.095 30.180 ;
        RECT 110.430 27.940 110.860 29.745 ;
        RECT 111.745 27.740 127.940 29.950 ;
        RECT 128.855 29.685 129.085 29.745 ;
        RECT 128.785 28.005 129.155 29.685 ;
        RECT 128.855 27.945 129.085 28.005 ;
        RECT 130.055 27.740 146.250 29.950 ;
        RECT 147.085 27.740 147.515 29.745 ;
        RECT 110.845 27.510 147.515 27.740 ;
        RECT 147.655 26.150 148.085 30.390 ;
        RECT 110.430 25.650 152.710 26.150 ;
        RECT 109.860 24.725 147.565 25.225 ;
        RECT 151.810 24.470 152.710 25.650 ;
        RECT 116.895 22.985 128.855 23.215 ;
        RECT 129.185 22.985 141.145 23.215 ;
        RECT 116.615 22.765 116.845 22.825 ;
        RECT 78.460 17.200 79.255 17.490 ;
        RECT 76.535 16.535 77.155 16.600 ;
        RECT 76.215 16.305 77.215 16.535 ;
        RECT 76.535 16.240 77.155 16.305 ;
        RECT 77.420 15.910 77.650 16.255 ;
        RECT 75.780 14.515 77.650 15.910 ;
        RECT 75.780 13.030 76.010 14.515 ;
        RECT 76.275 14.245 76.890 14.310 ;
        RECT 77.420 14.295 77.650 14.515 ;
        RECT 76.215 14.015 77.215 14.245 ;
        RECT 76.275 13.950 76.890 14.015 ;
        RECT 76.540 13.630 77.155 13.695 ;
        RECT 76.215 13.400 77.215 13.630 ;
        RECT 76.540 13.335 77.155 13.400 ;
        RECT 77.420 13.030 77.650 13.350 ;
        RECT 72.280 11.435 73.280 11.665 ;
        RECT 75.780 11.635 77.650 13.030 ;
        RECT 72.340 11.370 72.640 11.435 ;
        RECT 72.920 11.370 73.220 11.435 ;
        RECT 75.780 11.365 76.010 11.635 ;
        RECT 76.275 11.340 76.890 11.405 ;
        RECT 77.420 11.390 77.650 11.635 ;
        RECT 76.215 11.110 77.215 11.340 ;
        RECT 76.275 11.045 76.890 11.110 ;
        RECT 78.480 10.805 79.235 17.200 ;
        RECT 116.375 17.095 116.905 22.765 ;
        RECT 116.615 16.825 116.845 17.095 ;
        RECT 120.135 16.695 125.560 22.985 ;
        RECT 128.905 18.640 129.135 22.825 ;
        RECT 128.845 17.045 129.205 18.640 ;
        RECT 128.905 16.825 129.135 17.045 ;
        RECT 132.655 16.695 138.090 22.985 ;
        RECT 141.195 22.765 141.425 22.825 ;
        RECT 141.135 17.160 141.665 22.765 ;
        RECT 141.195 16.825 141.425 17.160 ;
        RECT 116.925 16.665 128.845 16.695 ;
        RECT 129.195 16.665 141.135 16.695 ;
        RECT 116.895 16.435 128.855 16.665 ;
        RECT 129.185 16.435 141.145 16.665 ;
        RECT 116.925 16.410 128.845 16.435 ;
        RECT 129.195 16.410 141.135 16.435 ;
        RECT 116.975 15.730 130.290 16.125 ;
        RECT 109.960 15.230 112.940 15.285 ;
        RECT 109.950 15.000 112.950 15.230 ;
        RECT 109.560 13.955 109.790 14.950 ;
        RECT 113.110 14.045 113.405 14.950 ;
        RECT 127.740 14.195 141.085 14.640 ;
        RECT 113.050 13.955 113.410 14.045 ;
        RECT 109.560 10.970 113.410 13.955 ;
        RECT 116.900 13.840 128.840 13.870 ;
        RECT 129.190 13.840 141.130 13.865 ;
        RECT 116.890 13.610 128.850 13.840 ;
        RECT 129.180 13.610 141.140 13.840 ;
        RECT 116.900 13.585 128.840 13.610 ;
        RECT 116.610 13.390 116.840 13.450 ;
        RECT 109.560 9.990 109.790 10.970 ;
        RECT 113.050 10.050 113.410 10.970 ;
        RECT 113.110 9.990 113.405 10.050 ;
        RECT 109.950 9.710 112.950 9.940 ;
        RECT 115.845 7.685 116.900 13.390 ;
        RECT 116.610 7.450 116.840 7.685 ;
        RECT 120.110 7.295 125.545 13.585 ;
        RECT 129.190 13.580 141.130 13.610 ;
        RECT 128.900 13.235 129.130 13.450 ;
        RECT 128.840 11.640 129.200 13.235 ;
        RECT 128.900 7.450 129.130 11.640 ;
        RECT 108.820 6.690 111.705 7.220 ;
        RECT 116.890 7.035 128.850 7.295 ;
        RECT 129.190 7.290 131.690 7.300 ;
        RECT 132.610 7.290 138.045 13.580 ;
        RECT 141.190 13.390 141.420 13.450 ;
        RECT 141.125 8.030 141.985 13.390 ;
        RECT 141.190 7.450 141.420 8.030 ;
        RECT 129.180 7.060 141.140 7.290 ;
        RECT 129.190 7.040 131.690 7.060 ;
        RECT 108.830 5.540 143.620 6.045 ;
      LAYER met2 ;
        RECT 52.080 48.485 53.050 48.720 ;
        RECT 51.050 47.960 53.050 48.485 ;
        RECT 77.975 48.340 81.975 48.640 ;
        RECT 51.050 47.690 67.055 47.960 ;
        RECT 51.050 43.040 53.050 47.690 ;
        RECT 66.785 47.075 67.055 47.690 ;
        RECT 54.205 46.620 55.305 46.940 ;
        RECT 66.785 46.910 68.170 47.075 ;
        RECT 70.640 47.050 74.400 47.855 ;
        RECT 64.490 46.650 68.170 46.910 ;
        RECT 63.115 46.235 63.715 46.355 ;
        RECT 61.145 45.975 61.505 46.215 ;
        RECT 60.145 45.715 61.505 45.975 ;
        RECT 63.115 45.975 63.725 46.235 ;
        RECT 57.085 45.350 58.185 45.630 ;
        RECT 60.145 45.475 60.505 45.715 ;
        RECT 58.290 44.685 58.650 44.925 ;
        RECT 58.290 44.425 59.780 44.685 ;
        RECT 51.050 42.780 55.305 43.040 ;
        RECT 51.050 35.300 53.050 42.780 ;
        RECT 54.205 38.880 55.305 39.200 ;
        RECT 55.965 35.975 56.565 44.330 ;
        RECT 59.420 44.185 59.780 44.425 ;
        RECT 61.610 42.750 62.710 43.070 ;
        RECT 58.290 42.105 58.650 42.345 ;
        RECT 58.290 41.845 60.505 42.105 ;
        RECT 60.145 41.605 60.505 41.845 ;
        RECT 61.145 40.815 61.505 41.555 ;
        RECT 59.420 40.555 61.505 40.815 ;
        RECT 57.085 40.190 58.185 40.470 ;
        RECT 59.420 40.315 59.780 40.555 ;
        RECT 63.115 39.845 63.715 45.975 ;
        RECT 66.785 44.415 68.170 46.650 ;
        RECT 64.485 44.060 65.585 44.340 ;
        RECT 66.785 42.655 67.445 44.415 ;
        RECT 69.715 43.510 72.815 43.880 ;
        RECT 73.450 42.655 74.400 47.050 ;
        RECT 75.630 45.315 76.055 47.110 ;
        RECT 77.905 46.640 81.975 48.340 ;
        RECT 77.905 46.510 79.970 46.640 ;
        RECT 77.810 46.250 79.970 46.510 ;
        RECT 77.905 45.210 79.970 46.250 ;
        RECT 76.230 44.950 79.970 45.210 ;
        RECT 75.630 43.045 76.055 44.840 ;
        RECT 77.905 43.375 79.970 44.950 ;
        RECT 66.785 41.885 74.400 42.655 ;
        RECT 64.490 41.480 65.590 41.760 ;
        RECT 63.110 39.585 63.715 39.845 ;
        RECT 63.115 38.565 63.715 39.585 ;
        RECT 66.785 39.170 67.445 41.885 ;
        RECT 76.230 41.585 77.030 41.905 ;
        RECT 72.290 41.400 72.690 41.430 ;
        RECT 72.250 40.590 72.720 41.400 ;
        RECT 64.490 38.910 67.445 39.170 ;
        RECT 61.145 38.235 61.505 38.475 ;
        RECT 63.105 38.305 63.715 38.565 ;
        RECT 60.145 37.975 61.505 38.235 ;
        RECT 57.085 37.610 58.185 37.890 ;
        RECT 60.145 37.735 60.505 37.975 ;
        RECT 58.290 36.945 58.650 37.345 ;
        RECT 58.290 36.685 59.780 36.945 ;
        RECT 59.420 36.445 59.780 36.685 ;
        RECT 55.960 35.715 56.565 35.975 ;
        RECT 51.050 35.040 55.305 35.300 ;
        RECT 51.050 27.565 53.050 35.040 ;
        RECT 55.965 34.665 56.565 35.715 ;
        RECT 61.610 35.010 62.710 35.330 ;
        RECT 55.965 34.405 56.570 34.665 ;
        RECT 54.205 31.140 55.305 31.460 ;
        RECT 55.965 28.200 56.565 34.405 ;
        RECT 58.290 34.365 58.650 34.605 ;
        RECT 58.290 34.105 60.505 34.365 ;
        RECT 60.145 33.865 60.505 34.105 ;
        RECT 61.145 33.075 61.505 33.735 ;
        RECT 59.420 32.815 61.505 33.075 ;
        RECT 57.085 32.450 58.185 32.730 ;
        RECT 59.420 32.575 59.780 32.815 ;
        RECT 63.115 30.825 63.715 38.305 ;
        RECT 64.490 36.320 65.590 36.600 ;
        RECT 64.490 33.740 65.590 34.020 ;
        RECT 66.785 31.430 67.445 38.910 ;
        RECT 64.490 31.170 67.445 31.430 ;
        RECT 61.145 30.495 61.505 30.735 ;
        RECT 60.145 30.235 61.505 30.495 ;
        RECT 63.115 30.565 63.725 30.825 ;
        RECT 57.085 29.870 58.185 30.150 ;
        RECT 60.145 29.995 60.505 30.235 ;
        RECT 63.115 30.140 63.715 30.565 ;
        RECT 63.110 29.880 63.715 30.140 ;
        RECT 58.290 29.205 58.650 29.575 ;
        RECT 58.290 28.945 59.780 29.205 ;
        RECT 59.420 28.705 59.780 28.945 ;
        RECT 55.965 27.940 56.575 28.200 ;
        RECT 51.050 27.305 55.305 27.565 ;
        RECT 51.050 19.820 53.050 27.305 ;
        RECT 55.965 26.940 56.565 27.940 ;
        RECT 61.610 27.270 62.710 27.590 ;
        RECT 55.960 26.680 56.565 26.940 ;
        RECT 54.205 23.400 55.305 23.720 ;
        RECT 55.965 20.485 56.565 26.680 ;
        RECT 58.290 26.625 58.650 26.865 ;
        RECT 58.290 26.365 60.505 26.625 ;
        RECT 60.145 26.125 60.505 26.365 ;
        RECT 61.145 25.335 61.505 25.995 ;
        RECT 59.420 25.075 61.505 25.335 ;
        RECT 57.085 24.710 58.185 24.990 ;
        RECT 59.420 24.835 59.780 25.075 ;
        RECT 63.115 24.345 63.715 29.880 ;
        RECT 64.490 28.580 65.590 28.860 ;
        RECT 64.490 26.000 65.590 26.280 ;
        RECT 63.115 24.085 63.725 24.345 ;
        RECT 61.145 22.755 61.505 22.995 ;
        RECT 60.145 22.495 61.505 22.755 ;
        RECT 57.085 22.130 58.185 22.410 ;
        RECT 60.145 22.255 60.505 22.495 ;
        RECT 58.290 21.465 58.650 21.830 ;
        RECT 58.290 21.205 59.780 21.465 ;
        RECT 59.420 20.965 59.780 21.205 ;
        RECT 55.950 20.225 56.565 20.485 ;
        RECT 51.050 19.560 55.305 19.820 ;
        RECT 51.050 5.515 53.050 19.560 ;
        RECT 55.965 19.175 56.565 20.225 ;
        RECT 61.610 19.530 62.710 19.850 ;
        RECT 55.960 18.915 56.565 19.175 ;
        RECT 54.205 15.660 55.305 15.980 ;
        RECT 55.965 14.890 56.565 18.915 ;
        RECT 58.290 18.885 58.650 19.125 ;
        RECT 58.290 18.625 60.505 18.885 ;
        RECT 60.145 18.385 60.505 18.625 ;
        RECT 61.145 17.595 61.505 18.255 ;
        RECT 59.420 17.335 61.505 17.595 ;
        RECT 57.085 16.970 58.185 17.250 ;
        RECT 59.420 17.095 59.780 17.335 ;
        RECT 63.115 16.610 63.715 24.085 ;
        RECT 66.785 23.690 67.445 31.170 ;
        RECT 64.490 23.430 67.445 23.690 ;
        RECT 64.490 20.840 65.590 21.120 ;
        RECT 64.490 18.260 65.590 18.540 ;
        RECT 58.290 16.305 58.650 16.545 ;
        RECT 61.145 16.305 61.505 16.545 ;
        RECT 63.105 16.350 63.715 16.610 ;
        RECT 58.290 16.045 59.780 16.305 ;
        RECT 59.420 15.805 59.780 16.045 ;
        RECT 60.145 16.045 61.505 16.305 ;
        RECT 60.145 15.805 60.505 16.045 ;
        RECT 63.115 14.890 63.715 16.350 ;
        RECT 66.785 15.950 67.445 23.430 ;
        RECT 64.490 15.690 67.445 15.950 ;
        RECT 66.785 15.305 67.445 15.690 ;
        RECT 55.965 14.290 63.715 14.890 ;
        RECT 70.490 11.005 71.545 38.505 ;
        RECT 72.290 37.220 72.690 40.590 ;
        RECT 77.895 40.585 79.970 43.375 ;
        RECT 76.410 40.325 79.970 40.585 ;
        RECT 76.230 39.005 77.030 39.325 ;
        RECT 77.895 38.445 79.970 40.325 ;
        RECT 78.635 36.755 79.970 38.445 ;
        RECT 72.290 30.770 72.690 36.190 ;
        RECT 78.460 35.900 79.970 36.755 ;
        RECT 76.490 35.640 79.970 35.900 ;
        RECT 72.870 33.610 73.270 34.900 ;
        RECT 72.870 33.350 76.890 33.610 ;
        RECT 72.870 32.060 73.270 33.350 ;
        RECT 72.290 24.320 72.690 29.740 ;
        RECT 78.460 29.450 79.970 35.640 ;
        RECT 108.350 33.885 154.395 35.880 ;
        RECT 108.350 33.880 151.230 33.885 ;
        RECT 76.490 29.190 79.970 29.450 ;
        RECT 72.870 27.160 73.270 28.450 ;
        RECT 72.870 26.900 76.890 27.160 ;
        RECT 72.870 25.610 73.270 26.900 ;
        RECT 72.290 17.870 72.690 23.290 ;
        RECT 78.460 23.000 79.970 29.190 ;
        RECT 110.380 26.165 110.810 29.745 ;
        RECT 128.835 27.955 129.105 33.880 ;
        RECT 110.380 25.645 111.975 26.165 ;
        RECT 114.470 25.650 116.275 26.150 ;
        RECT 139.790 25.650 141.615 26.150 ;
        RECT 76.490 22.740 79.970 23.000 ;
        RECT 72.870 20.710 73.270 22.000 ;
        RECT 72.870 20.450 76.890 20.710 ;
        RECT 72.870 19.160 73.270 20.450 ;
        RECT 78.460 17.625 79.970 22.740 ;
        RECT 72.290 11.680 72.690 16.840 ;
        RECT 78.430 16.550 79.970 17.625 ;
        RECT 76.485 16.290 79.970 16.550 ;
        RECT 72.870 14.260 73.270 15.550 ;
        RECT 72.870 14.000 76.935 14.260 ;
        RECT 72.870 12.710 73.270 14.000 ;
        RECT 78.430 13.645 79.970 16.290 ;
        RECT 110.010 14.960 112.890 15.385 ;
        RECT 113.100 14.090 113.360 14.095 ;
        RECT 76.490 13.385 79.970 13.645 ;
        RECT 72.290 11.420 75.420 11.680 ;
        RECT 74.530 11.355 75.420 11.420 ;
        RECT 74.530 11.095 76.940 11.355 ;
        RECT 74.530 9.060 75.420 11.095 ;
        RECT 78.430 9.895 79.970 13.385 ;
        RECT 113.085 10.000 113.375 14.090 ;
        RECT 115.845 13.440 116.275 25.650 ;
        RECT 116.425 24.725 118.355 25.225 ;
        RECT 116.425 19.875 116.855 24.725 ;
        RECT 141.185 19.875 141.615 25.650 ;
        RECT 147.135 25.225 147.565 29.745 ;
        RECT 141.765 24.725 143.635 25.225 ;
        RECT 145.460 24.725 147.565 25.225 ;
        RECT 128.875 16.945 129.155 18.755 ;
        RECT 116.975 15.770 118.025 16.745 ;
        RECT 127.740 13.535 128.790 14.580 ;
        RECT 129.240 13.530 130.290 16.185 ;
        RECT 140.035 14.205 141.085 16.745 ;
        RECT 141.765 13.440 142.195 24.725 ;
        RECT 151.860 24.420 152.660 26.150 ;
        RECT 115.845 10.570 116.850 13.440 ;
        RECT 128.870 11.540 129.160 13.335 ;
        RECT 74.720 9.015 75.205 9.060 ;
        RECT 115.845 7.685 116.860 10.570 ;
        RECT 141.175 7.980 142.195 13.440 ;
        RECT 108.340 7.515 112.250 7.520 ;
        RECT 66.720 6.065 112.250 7.515 ;
        RECT 116.950 6.970 119.350 7.360 ;
        RECT 129.240 6.980 131.640 7.370 ;
        RECT 66.720 5.520 143.560 6.065 ;
        RECT 66.720 5.515 89.070 5.520 ;
      LAYER met3 ;
        RECT 57.780 47.260 65.565 47.630 ;
        RECT 54.230 46.570 55.280 46.990 ;
        RECT 57.780 45.680 58.150 47.260 ;
        RECT 57.110 45.300 58.160 45.680 ;
        RECT 57.780 40.520 58.150 45.300 ;
        RECT 65.185 44.390 65.565 47.260 ;
        RECT 75.655 45.265 76.030 47.160 ;
        RECT 80.050 46.755 81.935 48.525 ;
        RECT 64.510 44.010 65.565 44.390 ;
        RECT 61.635 42.700 62.685 43.120 ;
        RECT 65.185 41.810 65.565 44.010 ;
        RECT 69.740 43.460 72.790 43.930 ;
        RECT 75.655 42.995 76.030 44.890 ;
        RECT 64.515 41.430 65.565 41.810 ;
        RECT 76.255 41.535 77.005 41.955 ;
        RECT 72.275 41.430 72.695 41.450 ;
        RECT 65.185 41.050 72.695 41.430 ;
        RECT 57.110 40.140 58.160 40.520 ;
        RECT 54.230 38.830 55.280 39.250 ;
        RECT 57.780 37.940 58.150 40.140 ;
        RECT 57.110 37.560 58.160 37.940 ;
        RECT 57.780 32.780 58.150 37.560 ;
        RECT 65.185 36.650 65.565 41.050 ;
        RECT 72.275 40.540 72.695 41.050 ;
        RECT 76.255 38.955 77.005 39.375 ;
        RECT 64.515 36.270 65.565 36.650 ;
        RECT 61.635 34.960 62.685 35.380 ;
        RECT 65.185 34.070 65.565 36.270 ;
        RECT 64.515 33.690 65.565 34.070 ;
        RECT 150.435 33.885 154.430 35.875 ;
        RECT 57.110 32.400 58.160 32.780 ;
        RECT 54.230 31.090 55.280 31.510 ;
        RECT 57.780 30.200 58.150 32.400 ;
        RECT 57.110 29.820 58.160 30.200 ;
        RECT 57.780 25.040 58.150 29.820 ;
        RECT 65.185 28.910 65.565 33.690 ;
        RECT 64.515 28.530 65.565 28.910 ;
        RECT 61.635 27.220 62.685 27.640 ;
        RECT 65.185 26.330 65.565 28.530 ;
        RECT 64.515 25.950 65.565 26.330 ;
        RECT 57.110 24.660 58.160 25.040 ;
        RECT 54.230 23.350 55.280 23.770 ;
        RECT 57.780 22.460 58.150 24.660 ;
        RECT 57.110 22.080 58.160 22.460 ;
        RECT 57.780 17.620 58.150 22.080 ;
        RECT 65.185 21.170 65.565 25.950 ;
        RECT 151.810 24.445 152.710 26.125 ;
        RECT 64.515 20.790 65.565 21.170 ;
        RECT 61.635 19.480 62.685 19.900 ;
        RECT 65.185 18.590 65.565 20.790 ;
        RECT 64.515 18.210 65.565 18.590 ;
        RECT 57.780 17.300 58.160 17.620 ;
        RECT 57.110 16.920 58.160 17.300 ;
        RECT 54.230 15.610 55.280 16.030 ;
        RECT 128.820 15.360 129.210 18.730 ;
        RECT 109.960 14.985 129.210 15.360 ;
        RECT 74.670 9.040 75.255 9.990 ;
        RECT 51.205 5.685 52.910 7.430 ;
        RECT 66.670 5.520 70.465 7.510 ;
        RECT 113.035 5.140 113.935 14.065 ;
        RECT 128.820 11.565 129.210 14.985 ;
        RECT 93.850 4.240 113.935 5.140 ;
        RECT 116.900 6.995 119.400 7.335 ;
        RECT 129.190 7.005 131.690 7.345 ;
        RECT 116.900 3.910 117.800 6.995 ;
        RECT 115.160 3.020 117.800 3.910 ;
        RECT 116.900 3.015 117.800 3.020 ;
        RECT 129.190 3.910 130.090 7.005 ;
        RECT 129.190 3.020 131.870 3.910 ;
        RECT 129.190 3.015 130.090 3.020 ;
      LAYER met4 ;
        RECT 30.670 220.760 30.970 224.760 ;
        RECT 33.430 220.760 33.730 224.760 ;
        RECT 36.190 220.760 36.490 224.760 ;
        RECT 38.950 220.760 39.250 224.760 ;
        RECT 41.710 220.760 42.010 224.760 ;
        RECT 44.470 220.760 44.770 224.760 ;
        RECT 47.230 220.760 47.530 224.760 ;
        RECT 49.990 220.760 50.290 224.760 ;
        RECT 52.750 220.760 53.050 224.760 ;
        RECT 55.510 220.760 55.810 224.760 ;
        RECT 58.270 220.760 58.570 224.760 ;
        RECT 61.030 220.760 61.330 224.760 ;
        RECT 63.790 220.760 64.090 224.760 ;
        RECT 66.550 220.760 66.850 224.760 ;
        RECT 69.310 220.760 69.610 224.760 ;
        RECT 72.070 220.760 72.370 224.760 ;
        RECT 74.830 220.760 75.130 224.760 ;
        RECT 77.590 220.760 77.890 224.760 ;
        RECT 80.350 220.760 80.650 224.760 ;
        RECT 83.110 220.760 83.410 224.760 ;
        RECT 85.870 220.760 86.170 224.760 ;
        RECT 88.630 220.760 88.930 224.760 ;
        RECT 91.390 220.760 91.690 224.760 ;
        RECT 94.150 220.760 94.450 224.760 ;
        RECT 4.000 218.760 94.450 220.760 ;
        RECT 57.905 48.920 76.020 49.300 ;
        RECT 57.905 48.360 58.290 48.920 ;
        RECT 54.250 47.980 62.035 48.360 ;
        RECT 54.250 46.945 54.630 47.980 ;
        RECT 54.250 46.615 55.260 46.945 ;
        RECT 54.250 39.205 54.630 46.615 ;
        RECT 61.655 43.075 62.035 47.980 ;
        RECT 69.760 43.505 72.790 43.885 ;
        RECT 61.655 42.745 62.665 43.075 ;
        RECT 54.250 38.875 55.260 39.205 ;
        RECT 54.250 31.465 54.630 38.875 ;
        RECT 61.655 35.335 62.035 42.745 ;
        RECT 72.410 40.605 72.790 43.505 ;
        RECT 75.655 42.855 76.020 48.920 ;
        RECT 79.975 46.640 157.000 48.640 ;
        RECT 74.750 41.580 76.985 41.910 ;
        RECT 74.750 40.605 75.130 41.580 ;
        RECT 72.410 40.275 75.130 40.605 ;
        RECT 74.750 39.330 75.130 40.275 ;
        RECT 74.750 39.000 76.985 39.330 ;
        RECT 61.655 35.005 62.665 35.335 ;
        RECT 54.250 31.135 55.260 31.465 ;
        RECT 54.250 23.725 54.630 31.135 ;
        RECT 61.655 27.595 62.035 35.005 ;
        RECT 150.025 33.880 157.000 35.880 ;
        RECT 61.655 27.265 62.665 27.595 ;
        RECT 54.250 23.395 55.260 23.725 ;
        RECT 54.250 15.985 54.630 23.395 ;
        RECT 61.655 19.855 62.035 27.265 ;
        RECT 61.655 19.525 62.665 19.855 ;
        RECT 54.250 15.655 55.260 15.985 ;
        RECT 74.715 9.960 75.210 9.970 ;
        RECT 4.000 5.515 70.420 7.515 ;
        RECT 74.530 1.000 75.430 9.960 ;
        RECT 93.850 4.240 96.385 5.140 ;
        RECT 93.850 1.000 94.750 4.240 ;
        RECT 113.170 3.015 117.800 3.915 ;
        RECT 129.190 3.015 133.390 3.915 ;
        RECT 113.170 1.000 114.070 3.015 ;
        RECT 132.490 1.000 133.390 3.015 ;
        RECT 151.810 1.000 152.710 26.150 ;
  END
END tt_um_DalinEM_diff_amp
END LIBRARY

