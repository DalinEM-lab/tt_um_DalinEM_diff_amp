magic
tech sky130A
magscale 1 2
timestamp 1740447052
<< nwell >>
rect -1003 -919 1003 919
<< pmos >>
rect -807 -700 -447 700
rect -389 -700 -29 700
rect 29 -700 389 700
rect 447 -700 807 700
<< pdiff >>
rect -865 688 -807 700
rect -865 -688 -853 688
rect -819 -688 -807 688
rect -865 -700 -807 -688
rect -447 688 -389 700
rect -447 -688 -435 688
rect -401 -688 -389 688
rect -447 -700 -389 -688
rect -29 688 29 700
rect -29 -688 -17 688
rect 17 -688 29 688
rect -29 -700 29 -688
rect 389 688 447 700
rect 389 -688 401 688
rect 435 -688 447 688
rect 389 -700 447 -688
rect 807 688 865 700
rect 807 -688 819 688
rect 853 -688 865 688
rect 807 -700 865 -688
<< pdiffc >>
rect -853 -688 -819 688
rect -435 -688 -401 688
rect -17 -688 17 688
rect 401 -688 435 688
rect 819 -688 853 688
<< nsubdiff >>
rect -967 849 -871 883
rect 871 849 967 883
rect -967 787 -933 849
rect 933 787 967 849
rect -967 -849 -933 -787
rect 933 -849 967 -787
rect -967 -883 -871 -849
rect 871 -883 967 -849
<< nsubdiffcont >>
rect -871 849 871 883
rect -967 -787 -933 787
rect 933 -787 967 787
rect -871 -883 871 -849
<< poly >>
rect -807 781 -447 797
rect -807 747 -791 781
rect -463 747 -447 781
rect -807 700 -447 747
rect -389 781 -29 797
rect -389 747 -373 781
rect -45 747 -29 781
rect -389 700 -29 747
rect 29 781 389 797
rect 29 747 45 781
rect 373 747 389 781
rect 29 700 389 747
rect 447 781 807 797
rect 447 747 463 781
rect 791 747 807 781
rect 447 700 807 747
rect -807 -747 -447 -700
rect -807 -781 -791 -747
rect -463 -781 -447 -747
rect -807 -797 -447 -781
rect -389 -747 -29 -700
rect -389 -781 -373 -747
rect -45 -781 -29 -747
rect -389 -797 -29 -781
rect 29 -747 389 -700
rect 29 -781 45 -747
rect 373 -781 389 -747
rect 29 -797 389 -781
rect 447 -747 807 -700
rect 447 -781 463 -747
rect 791 -781 807 -747
rect 447 -797 807 -781
<< polycont >>
rect -791 747 -463 781
rect -373 747 -45 781
rect 45 747 373 781
rect 463 747 791 781
rect -791 -781 -463 -747
rect -373 -781 -45 -747
rect 45 -781 373 -747
rect 463 -781 791 -747
<< locali >>
rect -967 849 -871 883
rect 871 849 967 883
rect -967 787 -933 849
rect 933 787 967 849
rect -807 747 -791 781
rect -463 747 -447 781
rect -389 747 -373 781
rect -45 747 -29 781
rect 29 747 45 781
rect 373 747 389 781
rect 447 747 463 781
rect 791 747 807 781
rect -853 688 -819 704
rect -853 -704 -819 -688
rect -435 688 -401 704
rect -435 -704 -401 -688
rect -17 688 17 704
rect -17 -704 17 -688
rect 401 688 435 704
rect 401 -704 435 -688
rect 819 688 853 704
rect 819 -704 853 -688
rect -807 -781 -791 -747
rect -463 -781 -447 -747
rect -389 -781 -373 -747
rect -45 -781 -29 -747
rect 29 -781 45 -747
rect 373 -781 389 -747
rect 447 -781 463 -747
rect 791 -781 807 -747
rect -967 -849 -933 -787
rect 933 -849 967 -787
rect -967 -883 -871 -849
rect 871 -883 967 -849
<< viali >>
rect -791 747 -463 781
rect -373 747 -45 781
rect 45 747 373 781
rect 463 747 791 781
rect -853 -688 -819 688
rect -435 -688 -401 688
rect -17 -688 17 688
rect 401 -688 435 688
rect 819 -688 853 688
rect -791 -781 -463 -747
rect -373 -781 -45 -747
rect 45 -781 373 -747
rect 463 -781 791 -747
<< metal1 >>
rect -803 781 -451 787
rect -803 747 -791 781
rect -463 747 -451 781
rect -803 741 -451 747
rect -385 781 -33 787
rect -385 747 -373 781
rect -45 747 -33 781
rect -385 741 -33 747
rect 33 781 385 787
rect 33 747 45 781
rect 373 747 385 781
rect 33 741 385 747
rect 451 781 803 787
rect 451 747 463 781
rect 791 747 803 781
rect 451 741 803 747
rect -859 688 -813 700
rect -859 -688 -853 688
rect -819 -688 -813 688
rect -859 -700 -813 -688
rect -441 688 -395 700
rect -441 -688 -435 688
rect -401 -688 -395 688
rect -441 -700 -395 -688
rect -23 688 23 700
rect -23 -688 -17 688
rect 17 -688 23 688
rect -23 -700 23 -688
rect 395 688 441 700
rect 395 -688 401 688
rect 435 -688 441 688
rect 395 -700 441 -688
rect 813 688 859 700
rect 813 -688 819 688
rect 853 -688 859 688
rect 813 -700 859 -688
rect -803 -747 -451 -741
rect -803 -781 -791 -747
rect -463 -781 -451 -747
rect -803 -787 -451 -781
rect -385 -747 -33 -741
rect -385 -781 -373 -747
rect -45 -781 -33 -747
rect -385 -787 -33 -781
rect 33 -747 385 -741
rect 33 -781 45 -747
rect 373 -781 385 -747
rect 33 -787 385 -781
rect 451 -747 803 -741
rect 451 -781 463 -747
rect 791 -781 803 -747
rect 451 -787 803 -781
<< properties >>
string FIXED_BBOX -950 -866 950 866
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.0 l 1.8 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
