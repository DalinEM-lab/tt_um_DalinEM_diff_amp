MACRO BGR_BJT_final
  CLASS BLOCK ;
  FOREIGN BGR_BJT_final ;
  ORIGIN 0.840 0.010 ;
  SIZE 39.405 BY 28.420 ;
  PIN vcc
    ANTENNADIFFAREA 17.077549 ;
    PORT
      LAYER met2 ;
        RECT 38.550 0.960 38.560 0.970 ;
    END
  END vcc
  PIN vss
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 55.184998 ;
    PORT
      LAYER met2 ;
        RECT -0.260 27.565 -0.250 27.575 ;
    END
  END vss
  PIN vref
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met2 ;
        RECT 38.325 5.185 38.335 5.195 ;
    END
  END vref
  OBS
      LAYER pwell ;
        RECT -0.005 21.815 34.205 28.035 ;
        RECT -0.005 21.795 10.795 21.815 ;
        RECT 10.955 21.795 34.205 21.815 ;
        RECT -0.005 21.565 34.205 21.795 ;
        RECT -0.005 21.550 10.785 21.565 ;
        RECT 10.950 21.550 34.205 21.565 ;
        RECT -0.005 12.465 34.205 21.550 ;
        RECT 0.265 11.470 6.965 12.235 ;
        RECT 0.265 6.300 1.030 11.470 ;
        RECT 6.200 6.300 6.965 11.470 ;
        RECT 0.265 5.535 6.965 6.300 ;
        RECT 9.800 5.255 38.170 9.490 ;
      LAYER nwell ;
        RECT 0.065 4.990 5.985 4.995 ;
        RECT 0.065 1.835 10.140 4.990 ;
        RECT 11.855 1.840 15.815 5.030 ;
        RECT 18.305 1.840 22.265 5.030 ;
        RECT 24.755 1.840 28.715 5.030 ;
        RECT 0.085 1.830 10.140 1.835 ;
        RECT 31.235 1.775 38.100 4.950 ;
      LAYER li1 ;
        RECT -0.030 26.605 33.560 28.410 ;
        RECT 0.405 13.540 0.865 26.605 ;
        RECT 1.825 26.145 2.825 26.315 ;
        RECT 3.115 26.145 4.115 26.315 ;
        RECT 4.405 26.145 5.405 26.315 ;
        RECT 5.695 26.145 6.695 26.315 ;
        RECT 6.985 26.145 7.985 26.315 ;
        RECT 8.275 26.145 9.275 26.315 ;
        RECT 9.565 26.145 10.565 26.315 ;
        RECT 10.855 26.145 11.855 26.315 ;
        RECT 12.145 26.145 13.145 26.315 ;
        RECT 13.435 26.145 14.435 26.315 ;
        RECT 14.725 26.145 15.725 26.315 ;
        RECT 16.015 26.145 17.015 26.315 ;
        RECT 17.305 26.145 18.305 26.315 ;
        RECT 18.595 26.145 19.595 26.315 ;
        RECT 19.885 26.145 20.885 26.315 ;
        RECT 21.175 26.145 22.175 26.315 ;
        RECT 22.465 26.145 23.465 26.315 ;
        RECT 23.755 26.145 24.755 26.315 ;
        RECT 25.045 26.145 26.045 26.315 ;
        RECT 26.335 26.145 27.335 26.315 ;
        RECT 27.625 26.145 28.625 26.315 ;
        RECT 28.915 26.145 29.915 26.315 ;
        RECT 30.205 26.145 31.205 26.315 ;
        RECT 31.495 26.145 32.495 26.315 ;
        RECT 1.595 21.935 1.765 25.975 ;
        RECT 2.885 21.935 3.055 25.975 ;
        RECT 4.175 21.935 4.345 25.975 ;
        RECT 5.465 21.935 5.635 25.975 ;
        RECT 6.755 21.935 6.925 25.975 ;
        RECT 8.045 21.935 8.215 25.975 ;
        RECT 9.335 21.935 9.505 25.975 ;
        RECT 10.625 21.935 10.795 25.975 ;
        RECT 11.915 21.935 12.085 25.975 ;
        RECT 13.205 21.935 13.375 25.975 ;
        RECT 14.495 21.935 14.665 25.975 ;
        RECT 15.785 21.935 15.955 25.975 ;
        RECT 17.075 21.935 17.245 25.975 ;
        RECT 18.365 21.935 18.535 25.975 ;
        RECT 19.655 21.935 19.825 25.975 ;
        RECT 20.945 21.935 21.115 25.975 ;
        RECT 22.235 21.935 22.405 25.975 ;
        RECT 23.525 21.935 23.695 25.975 ;
        RECT 24.815 21.935 24.985 25.975 ;
        RECT 26.105 21.935 26.275 25.975 ;
        RECT 27.395 21.935 27.565 25.975 ;
        RECT 28.685 21.935 28.855 25.975 ;
        RECT 29.975 21.935 30.145 25.975 ;
        RECT 31.265 21.935 31.435 25.975 ;
        RECT 32.555 21.935 32.725 25.975 ;
        RECT 1.825 21.595 2.825 21.765 ;
        RECT 3.115 21.595 4.115 21.765 ;
        RECT 4.405 21.595 5.405 21.765 ;
        RECT 5.695 21.595 6.695 21.765 ;
        RECT 6.985 21.595 7.985 21.765 ;
        RECT 8.275 21.595 9.275 21.765 ;
        RECT 9.565 21.595 10.565 21.765 ;
        RECT 10.855 21.595 11.855 21.765 ;
        RECT 12.145 21.595 13.145 21.765 ;
        RECT 13.435 21.595 14.435 21.765 ;
        RECT 14.725 21.595 15.725 21.765 ;
        RECT 16.015 21.595 17.015 21.765 ;
        RECT 17.305 21.595 18.305 21.765 ;
        RECT 18.595 21.595 19.595 21.765 ;
        RECT 19.885 21.595 20.885 21.765 ;
        RECT 21.175 21.595 22.175 21.765 ;
        RECT 22.465 21.595 23.465 21.765 ;
        RECT 23.755 21.595 24.755 21.765 ;
        RECT 25.045 21.595 26.045 21.765 ;
        RECT 26.335 21.595 27.335 21.765 ;
        RECT 27.625 21.595 28.625 21.765 ;
        RECT 28.915 21.595 29.915 21.765 ;
        RECT 30.205 21.595 31.205 21.765 ;
        RECT 31.495 21.595 32.495 21.765 ;
        RECT 1.825 18.740 2.825 18.910 ;
        RECT 3.115 18.740 4.115 18.910 ;
        RECT 4.405 18.740 5.405 18.910 ;
        RECT 5.695 18.740 6.695 18.910 ;
        RECT 6.985 18.740 7.985 18.910 ;
        RECT 8.275 18.740 9.275 18.910 ;
        RECT 9.565 18.740 10.565 18.910 ;
        RECT 10.855 18.740 11.855 18.910 ;
        RECT 12.145 18.740 13.145 18.910 ;
        RECT 13.435 18.740 14.435 18.910 ;
        RECT 14.725 18.740 15.725 18.910 ;
        RECT 16.015 18.740 17.015 18.910 ;
        RECT 17.305 18.740 18.305 18.910 ;
        RECT 18.595 18.740 19.595 18.910 ;
        RECT 19.885 18.740 20.885 18.910 ;
        RECT 21.175 18.740 22.175 18.910 ;
        RECT 22.465 18.740 23.465 18.910 ;
        RECT 23.755 18.740 24.755 18.910 ;
        RECT 25.045 18.740 26.045 18.910 ;
        RECT 26.335 18.740 27.335 18.910 ;
        RECT 27.625 18.740 28.625 18.910 ;
        RECT 28.915 18.740 29.915 18.910 ;
        RECT 30.205 18.740 31.205 18.910 ;
        RECT 31.495 18.740 32.495 18.910 ;
        RECT 1.595 14.530 1.765 18.570 ;
        RECT 2.885 14.530 3.055 18.570 ;
        RECT 4.175 14.530 4.345 18.570 ;
        RECT 5.465 14.530 5.635 18.570 ;
        RECT 6.755 14.530 6.925 18.570 ;
        RECT 8.045 14.530 8.215 18.570 ;
        RECT 9.335 14.530 9.505 18.570 ;
        RECT 10.625 14.530 10.795 18.570 ;
        RECT 11.915 14.530 12.085 18.570 ;
        RECT 13.205 14.530 13.375 18.570 ;
        RECT 14.495 14.530 14.665 18.570 ;
        RECT 15.785 14.530 15.955 18.570 ;
        RECT 17.075 14.530 17.245 18.570 ;
        RECT 18.365 14.530 18.535 18.570 ;
        RECT 19.655 14.530 19.825 18.570 ;
        RECT 20.945 14.530 21.115 18.570 ;
        RECT 22.235 14.530 22.405 18.570 ;
        RECT 23.525 14.530 23.695 18.570 ;
        RECT 24.815 14.530 24.985 18.570 ;
        RECT 26.105 14.530 26.275 18.570 ;
        RECT 27.395 14.530 27.565 18.570 ;
        RECT 28.685 14.530 28.855 18.570 ;
        RECT 29.975 14.530 30.145 18.570 ;
        RECT 31.265 14.530 31.435 18.570 ;
        RECT 32.555 14.530 32.725 18.570 ;
        RECT 1.825 14.190 2.825 14.360 ;
        RECT 3.115 14.190 4.115 14.360 ;
        RECT 4.405 14.190 5.405 14.360 ;
        RECT 5.695 14.190 6.695 14.360 ;
        RECT 6.985 14.190 7.985 14.360 ;
        RECT 8.275 14.190 9.275 14.360 ;
        RECT 9.565 14.190 10.565 14.360 ;
        RECT 10.855 14.190 11.855 14.360 ;
        RECT 12.145 14.190 13.145 14.360 ;
        RECT 13.435 14.190 14.435 14.360 ;
        RECT 14.725 14.190 15.725 14.360 ;
        RECT 16.015 14.190 17.015 14.360 ;
        RECT 17.305 14.190 18.305 14.360 ;
        RECT 18.595 14.190 19.595 14.360 ;
        RECT 19.885 14.190 20.885 14.360 ;
        RECT 21.175 14.190 22.175 14.360 ;
        RECT 22.465 14.190 23.465 14.360 ;
        RECT 23.755 14.190 24.755 14.360 ;
        RECT 25.045 14.190 26.045 14.360 ;
        RECT 26.335 14.190 27.335 14.360 ;
        RECT 27.625 14.190 28.625 14.360 ;
        RECT 28.915 14.190 29.915 14.360 ;
        RECT 30.205 14.190 31.205 14.360 ;
        RECT 31.495 14.190 32.495 14.360 ;
        RECT 32.980 13.575 33.560 26.605 ;
        RECT 1.665 13.540 33.560 13.575 ;
        RECT 0.405 12.535 33.560 13.540 ;
        RECT 0.400 12.105 33.560 12.535 ;
        RECT 0.395 12.075 33.560 12.105 ;
        RECT 0.395 10.930 6.835 12.075 ;
        RECT 0.395 6.840 1.570 10.930 ;
        RECT 1.880 7.150 5.350 10.620 ;
        RECT 5.660 6.840 6.835 10.930 ;
        RECT 9.950 9.750 33.560 12.075 ;
        RECT 9.950 9.705 38.065 9.750 ;
        RECT 0.395 5.665 6.835 6.840 ;
        RECT 9.955 8.470 38.065 9.705 ;
        RECT 9.955 5.995 10.570 8.470 ;
        RECT 11.255 8.060 12.255 8.230 ;
        RECT 12.545 8.060 13.545 8.230 ;
        RECT 13.835 8.060 14.835 8.230 ;
        RECT 15.125 8.060 16.125 8.230 ;
        RECT 16.415 8.060 17.415 8.230 ;
        RECT 17.705 8.060 18.705 8.230 ;
        RECT 18.995 8.060 19.995 8.230 ;
        RECT 20.285 8.060 21.285 8.230 ;
        RECT 21.575 8.060 22.575 8.230 ;
        RECT 22.865 8.060 23.865 8.230 ;
        RECT 24.155 8.060 25.155 8.230 ;
        RECT 25.445 8.060 26.445 8.230 ;
        RECT 26.735 8.060 27.735 8.230 ;
        RECT 28.025 8.060 29.025 8.230 ;
        RECT 29.315 8.060 30.315 8.230 ;
        RECT 30.605 8.060 31.605 8.230 ;
        RECT 31.895 8.060 32.895 8.230 ;
        RECT 33.185 8.060 34.185 8.230 ;
        RECT 34.475 8.060 35.475 8.230 ;
        RECT 35.765 8.060 36.765 8.230 ;
        RECT 11.025 6.850 11.195 7.890 ;
        RECT 12.315 6.850 12.485 7.890 ;
        RECT 13.605 6.850 13.775 7.890 ;
        RECT 14.895 6.850 15.065 7.890 ;
        RECT 16.185 6.850 16.355 7.890 ;
        RECT 17.475 6.850 17.645 7.890 ;
        RECT 18.765 6.850 18.935 7.890 ;
        RECT 20.055 6.850 20.225 7.890 ;
        RECT 21.345 6.850 21.515 7.890 ;
        RECT 22.635 6.850 22.805 7.890 ;
        RECT 23.925 6.850 24.095 7.890 ;
        RECT 25.215 6.850 25.385 7.890 ;
        RECT 26.505 6.850 26.675 7.890 ;
        RECT 27.795 6.850 27.965 7.890 ;
        RECT 29.085 6.850 29.255 7.890 ;
        RECT 30.375 6.850 30.545 7.890 ;
        RECT 31.665 6.850 31.835 7.890 ;
        RECT 32.955 6.850 33.125 7.890 ;
        RECT 34.245 6.850 34.415 7.890 ;
        RECT 35.535 6.850 35.705 7.890 ;
        RECT 36.825 6.850 36.995 7.890 ;
        RECT 11.255 6.510 12.255 6.680 ;
        RECT 12.545 6.510 13.545 6.680 ;
        RECT 13.835 6.510 14.835 6.680 ;
        RECT 15.125 6.510 16.125 6.680 ;
        RECT 16.415 6.510 17.415 6.680 ;
        RECT 17.705 6.510 18.705 6.680 ;
        RECT 18.995 6.510 19.995 6.680 ;
        RECT 20.285 6.510 21.285 6.680 ;
        RECT 21.575 6.510 22.575 6.680 ;
        RECT 22.865 6.510 23.865 6.680 ;
        RECT 24.155 6.510 25.155 6.680 ;
        RECT 25.445 6.510 26.445 6.680 ;
        RECT 26.735 6.510 27.735 6.680 ;
        RECT 28.025 6.510 29.025 6.680 ;
        RECT 29.315 6.510 30.315 6.680 ;
        RECT 30.605 6.510 31.605 6.680 ;
        RECT 31.895 6.510 32.895 6.680 ;
        RECT 33.185 6.510 34.185 6.680 ;
        RECT 34.475 6.510 35.475 6.680 ;
        RECT 35.765 6.510 36.765 6.680 ;
        RECT 37.450 5.995 38.065 8.470 ;
        RECT 9.955 5.300 38.065 5.995 ;
        RECT 11.930 4.950 15.765 4.960 ;
        RECT 0.255 4.560 9.960 4.800 ;
        RECT 0.255 2.340 0.515 4.560 ;
        RECT 1.235 4.165 3.235 4.335 ;
        RECT 3.525 4.165 5.525 4.335 ;
        RECT 6.860 4.165 7.860 4.335 ;
        RECT 8.150 4.165 9.150 4.335 ;
        RECT 1.005 3.410 1.175 3.950 ;
        RECT 3.295 3.410 3.465 3.950 ;
        RECT 5.585 3.410 5.755 3.950 ;
        RECT 1.235 3.025 3.235 3.195 ;
        RECT 3.525 3.025 5.525 3.195 ;
        RECT 6.630 2.910 6.800 3.950 ;
        RECT 7.920 2.910 8.090 3.950 ;
        RECT 9.210 2.910 9.380 3.950 ;
        RECT 6.860 2.525 7.860 2.695 ;
        RECT 8.150 2.525 9.150 2.695 ;
        RECT 9.715 2.655 9.960 4.560 ;
        RECT 11.920 4.620 15.765 4.950 ;
        RECT 11.920 2.655 12.310 4.620 ;
        RECT 12.835 4.170 14.835 4.340 ;
        RECT 15.370 4.040 15.760 4.620 ;
        RECT 18.315 4.550 22.265 4.930 ;
        RECT 18.335 4.040 18.760 4.550 ;
        RECT 19.285 4.170 21.285 4.340 ;
        RECT 12.605 2.915 12.775 3.955 ;
        RECT 14.895 2.915 15.065 3.955 ;
        RECT -0.130 2.335 1.070 2.340 ;
        RECT 1.300 2.335 6.240 2.340 ;
        RECT -0.130 2.325 6.240 2.335 ;
        RECT 9.555 2.325 12.325 2.655 ;
        RECT 12.835 2.530 14.835 2.700 ;
        RECT -0.130 2.290 12.325 2.325 ;
        RECT 15.370 2.290 18.760 4.040 ;
        RECT 21.865 4.100 22.265 4.550 ;
        RECT 24.795 4.560 28.715 4.975 ;
        RECT 31.265 4.920 38.115 4.930 ;
        RECT 24.795 4.100 25.250 4.560 ;
        RECT 25.735 4.170 27.735 4.340 ;
        RECT 19.055 2.915 19.225 3.955 ;
        RECT 21.345 2.915 21.515 3.955 ;
        RECT 19.285 2.530 21.285 2.700 ;
        RECT 21.865 2.295 25.250 4.100 ;
        RECT 28.235 4.100 28.715 4.560 ;
        RECT 31.255 4.535 38.115 4.920 ;
        RECT 31.255 4.100 31.680 4.535 ;
        RECT 32.185 4.170 34.185 4.340 ;
        RECT 35.090 4.170 37.090 4.340 ;
        RECT 25.505 2.915 25.675 3.955 ;
        RECT 27.795 2.915 27.965 3.955 ;
        RECT 25.735 2.530 27.735 2.700 ;
        RECT 28.235 2.295 31.680 4.100 ;
        RECT 31.955 2.915 32.125 3.955 ;
        RECT 34.245 2.915 34.415 3.955 ;
        RECT 34.860 2.915 35.030 3.955 ;
        RECT 37.150 2.915 37.320 3.955 ;
        RECT 32.185 2.530 34.185 2.700 ;
        RECT 35.090 2.530 37.090 2.700 ;
        RECT 21.865 2.290 25.730 2.295 ;
        RECT 28.230 2.290 31.680 2.295 ;
        RECT 37.595 2.290 38.115 4.535 ;
        RECT -0.130 2.210 38.115 2.290 ;
        RECT -0.130 0.790 38.110 2.210 ;
        RECT -0.130 0.170 38.145 0.790 ;
        RECT -0.125 0.000 38.145 0.170 ;
        RECT -0.125 -0.010 10.175 0.000 ;
      LAYER met1 ;
        RECT 0.425 27.120 33.435 28.050 ;
        RECT 0.470 26.740 0.800 26.800 ;
        RECT 0.450 25.980 0.820 26.740 ;
        RECT 1.845 26.115 4.095 26.345 ;
        RECT 4.425 26.115 6.675 26.345 ;
        RECT 7.005 26.115 11.835 26.345 ;
        RECT 12.165 26.115 14.415 26.345 ;
        RECT 14.745 26.115 19.575 26.345 ;
        RECT 19.905 26.115 22.155 26.345 ;
        RECT 22.485 26.115 27.315 26.345 ;
        RECT 27.645 26.115 29.895 26.345 ;
        RECT 30.225 26.115 32.475 26.345 ;
        RECT 0.470 25.920 0.800 25.980 ;
        RECT 1.565 25.895 1.795 25.955 ;
        RECT 1.470 24.895 1.890 25.895 ;
        RECT 1.565 21.955 1.795 24.895 ;
        RECT 0.470 21.790 0.800 21.850 ;
        RECT 2.090 21.795 2.535 26.115 ;
        RECT 2.855 23.015 3.085 25.955 ;
        RECT 2.780 22.015 3.160 23.015 ;
        RECT 2.855 21.955 3.085 22.015 ;
        RECT 3.410 21.810 3.855 26.115 ;
        RECT 4.145 24.135 4.375 25.955 ;
        RECT 4.080 23.635 4.440 24.135 ;
        RECT 4.145 21.955 4.375 23.635 ;
        RECT 3.410 21.795 4.085 21.810 ;
        RECT 4.655 21.795 5.100 26.115 ;
        RECT 5.435 25.895 5.665 25.955 ;
        RECT 5.370 24.895 5.730 25.895 ;
        RECT 5.435 21.955 5.665 24.895 ;
        RECT 5.975 21.810 6.415 26.115 ;
        RECT 6.725 24.135 6.955 25.955 ;
        RECT 6.660 23.635 7.020 24.135 ;
        RECT 6.725 21.955 6.955 23.635 ;
        RECT 5.975 21.795 6.665 21.810 ;
        RECT 7.280 21.795 7.720 26.115 ;
        RECT 8.015 23.015 8.245 25.955 ;
        RECT 7.940 22.015 8.320 23.015 ;
        RECT 8.015 21.955 8.245 22.015 ;
        RECT 8.595 21.795 9.035 26.115 ;
        RECT 9.305 25.895 9.535 25.955 ;
        RECT 9.210 24.895 9.630 25.895 ;
        RECT 9.305 21.955 9.535 24.895 ;
        RECT 9.845 21.795 10.285 26.115 ;
        RECT 10.595 23.015 10.825 25.955 ;
        RECT 10.520 22.015 10.900 23.015 ;
        RECT 10.595 21.955 10.825 22.015 ;
        RECT 11.140 21.860 11.580 26.115 ;
        RECT 11.885 24.135 12.115 25.955 ;
        RECT 11.820 23.635 12.180 24.135 ;
        RECT 11.885 21.955 12.115 23.635 ;
        RECT 11.030 21.810 11.580 21.860 ;
        RECT 11.030 21.795 11.825 21.810 ;
        RECT 12.405 21.795 12.870 26.115 ;
        RECT 13.175 25.895 13.405 25.955 ;
        RECT 13.110 24.895 13.470 25.895 ;
        RECT 13.175 21.955 13.405 24.895 ;
        RECT 13.715 21.810 14.155 26.115 ;
        RECT 14.465 24.135 14.695 25.955 ;
        RECT 14.400 23.635 14.760 24.135 ;
        RECT 14.465 21.955 14.695 23.635 ;
        RECT 13.715 21.795 14.405 21.810 ;
        RECT 15.040 21.795 15.480 26.115 ;
        RECT 15.755 23.015 15.985 25.955 ;
        RECT 15.680 22.015 16.060 23.015 ;
        RECT 15.755 21.955 15.985 22.015 ;
        RECT 16.320 21.795 16.760 26.115 ;
        RECT 17.045 25.895 17.275 25.955 ;
        RECT 16.950 24.895 17.370 25.895 ;
        RECT 17.045 21.955 17.275 24.895 ;
        RECT 17.605 21.795 18.045 26.115 ;
        RECT 18.335 23.015 18.565 25.955 ;
        RECT 18.260 22.015 18.640 23.015 ;
        RECT 18.335 21.955 18.565 22.015 ;
        RECT 18.900 21.810 19.340 26.115 ;
        RECT 19.625 24.135 19.855 25.955 ;
        RECT 19.560 23.635 19.920 24.135 ;
        RECT 19.625 21.955 19.855 23.635 ;
        RECT 18.815 21.795 19.565 21.810 ;
        RECT 20.160 21.795 20.600 26.115 ;
        RECT 20.915 25.895 21.145 25.955 ;
        RECT 20.845 24.895 21.205 25.895 ;
        RECT 20.915 21.955 21.145 24.895 ;
        RECT 21.445 21.810 21.885 26.115 ;
        RECT 22.205 24.135 22.435 25.955 ;
        RECT 22.140 23.635 22.500 24.135 ;
        RECT 22.205 21.955 22.435 23.635 ;
        RECT 21.445 21.795 22.145 21.810 ;
        RECT 22.780 21.795 23.220 26.115 ;
        RECT 23.495 23.015 23.725 25.955 ;
        RECT 23.420 22.015 23.800 23.015 ;
        RECT 23.495 21.955 23.725 22.015 ;
        RECT 24.000 21.795 24.440 26.115 ;
        RECT 24.785 25.895 25.015 25.955 ;
        RECT 24.690 24.895 25.110 25.895 ;
        RECT 24.785 21.955 25.015 24.895 ;
        RECT 25.325 21.795 25.765 26.115 ;
        RECT 26.075 23.015 26.305 25.955 ;
        RECT 26.000 22.015 26.380 23.015 ;
        RECT 26.075 21.955 26.305 22.015 ;
        RECT 26.580 21.810 27.020 26.115 ;
        RECT 27.365 24.135 27.595 25.955 ;
        RECT 27.300 23.635 27.660 24.135 ;
        RECT 27.365 21.955 27.595 23.635 ;
        RECT 26.580 21.795 27.305 21.810 ;
        RECT 27.910 21.795 28.350 26.115 ;
        RECT 28.655 25.895 28.885 25.955 ;
        RECT 28.590 24.895 28.950 25.895 ;
        RECT 28.655 21.955 28.885 24.895 ;
        RECT 29.195 21.810 29.635 26.115 ;
        RECT 29.945 24.135 30.175 25.955 ;
        RECT 29.880 23.635 30.240 24.135 ;
        RECT 29.945 21.955 30.175 23.635 ;
        RECT 29.195 21.795 29.885 21.810 ;
        RECT 30.565 21.795 31.005 26.115 ;
        RECT 31.235 23.015 31.465 25.955 ;
        RECT 31.160 22.015 31.540 23.015 ;
        RECT 31.235 21.955 31.465 22.015 ;
        RECT 31.780 21.810 32.220 26.115 ;
        RECT 32.525 25.895 32.755 25.955 ;
        RECT 32.430 24.895 32.850 25.895 ;
        RECT 32.525 21.955 32.755 24.895 ;
        RECT 31.780 21.795 32.465 21.810 ;
        RECT 0.450 21.050 0.820 21.790 ;
        RECT 1.845 21.565 4.095 21.795 ;
        RECT 4.425 21.565 6.675 21.795 ;
        RECT 7.005 21.565 11.835 21.795 ;
        RECT 12.165 21.565 14.415 21.795 ;
        RECT 14.745 21.565 19.575 21.795 ;
        RECT 19.905 21.565 22.155 21.795 ;
        RECT 22.485 21.565 27.315 21.795 ;
        RECT 27.645 21.565 29.895 21.795 ;
        RECT 30.225 21.565 32.475 21.795 ;
        RECT 3.485 21.550 4.085 21.565 ;
        RECT 6.065 21.550 6.665 21.565 ;
        RECT 11.030 21.550 11.825 21.565 ;
        RECT 13.805 21.550 14.405 21.565 ;
        RECT 18.815 21.550 19.565 21.565 ;
        RECT 21.545 21.550 22.145 21.565 ;
        RECT 26.600 21.550 27.305 21.565 ;
        RECT 29.285 21.550 29.885 21.565 ;
        RECT 31.865 21.550 32.465 21.565 ;
        RECT 11.030 21.500 11.255 21.550 ;
        RECT 0.470 20.990 0.800 21.050 ;
        RECT 0.920 20.420 32.705 20.680 ;
        RECT 0.920 10.410 1.180 20.420 ;
        RECT 1.875 19.695 32.705 19.955 ;
        RECT 2.195 18.940 2.795 18.955 ;
        RECT 6.855 18.940 7.955 18.955 ;
        RECT 9.935 18.940 10.535 18.955 ;
        RECT 14.675 18.940 15.695 18.955 ;
        RECT 17.675 18.940 18.275 18.955 ;
        RECT 22.415 18.940 23.435 18.955 ;
        RECT 25.415 18.940 26.015 18.955 ;
        RECT 30.155 18.940 31.175 18.955 ;
        RECT 31.865 18.940 32.465 18.955 ;
        RECT 1.845 18.710 2.805 18.940 ;
        RECT 3.135 18.710 7.965 18.940 ;
        RECT 8.295 18.710 10.545 18.940 ;
        RECT 10.875 18.710 15.705 18.940 ;
        RECT 16.035 18.710 18.285 18.940 ;
        RECT 18.615 18.710 23.445 18.940 ;
        RECT 23.775 18.710 26.025 18.940 ;
        RECT 26.355 18.710 31.185 18.940 ;
        RECT 31.515 18.710 32.475 18.940 ;
        RECT 2.130 18.695 2.795 18.710 ;
        RECT 1.565 15.610 1.795 18.550 ;
        RECT 1.500 14.610 1.860 15.610 ;
        RECT 1.565 14.550 1.795 14.610 ;
        RECT 2.130 14.390 2.570 18.695 ;
        RECT 2.855 16.985 3.085 18.550 ;
        RECT 2.790 16.485 3.150 16.985 ;
        RECT 2.855 14.550 3.085 16.485 ;
        RECT 3.390 14.390 3.830 18.710 ;
        RECT 4.145 15.615 4.375 18.550 ;
        RECT 4.070 14.615 4.450 15.615 ;
        RECT 4.145 14.550 4.375 14.615 ;
        RECT 4.635 14.390 5.075 18.710 ;
        RECT 5.435 18.490 5.665 18.550 ;
        RECT 5.340 17.490 5.760 18.490 ;
        RECT 5.435 14.550 5.665 17.490 ;
        RECT 5.985 14.390 6.425 18.710 ;
        RECT 6.855 18.695 7.955 18.710 ;
        RECT 6.725 15.610 6.955 18.550 ;
        RECT 6.650 14.610 7.030 15.610 ;
        RECT 6.725 14.550 6.955 14.610 ;
        RECT 7.230 14.390 7.670 18.695 ;
        RECT 8.015 16.985 8.245 18.550 ;
        RECT 7.950 16.485 8.310 16.985 ;
        RECT 8.015 14.550 8.245 16.485 ;
        RECT 8.545 14.390 8.985 18.710 ;
        RECT 9.815 18.695 10.535 18.710 ;
        RECT 9.305 15.610 9.535 18.550 ;
        RECT 9.240 14.610 9.600 15.610 ;
        RECT 9.305 14.550 9.535 14.610 ;
        RECT 9.815 14.390 10.255 18.695 ;
        RECT 10.595 16.985 10.825 18.550 ;
        RECT 10.530 16.485 10.890 16.985 ;
        RECT 10.595 14.550 10.825 16.485 ;
        RECT 11.150 14.390 11.590 18.710 ;
        RECT 11.885 15.610 12.115 18.550 ;
        RECT 11.810 14.610 12.190 15.610 ;
        RECT 11.885 14.550 12.115 14.610 ;
        RECT 12.415 14.390 12.855 18.710 ;
        RECT 13.175 18.490 13.405 18.550 ;
        RECT 13.080 17.490 13.500 18.490 ;
        RECT 13.175 14.550 13.405 17.490 ;
        RECT 13.675 14.390 14.115 18.710 ;
        RECT 14.675 18.695 15.695 18.710 ;
        RECT 14.465 15.610 14.695 18.550 ;
        RECT 14.390 14.610 14.770 15.610 ;
        RECT 14.465 14.550 14.695 14.610 ;
        RECT 15.030 14.390 15.470 18.695 ;
        RECT 15.755 16.985 15.985 18.550 ;
        RECT 15.690 16.485 16.050 16.985 ;
        RECT 15.755 14.550 15.985 16.485 ;
        RECT 16.260 14.390 16.665 18.710 ;
        RECT 17.560 18.695 18.275 18.710 ;
        RECT 17.045 15.610 17.275 18.550 ;
        RECT 16.980 14.610 17.340 15.610 ;
        RECT 17.045 14.550 17.275 14.610 ;
        RECT 17.560 14.390 17.965 18.695 ;
        RECT 18.335 16.990 18.565 18.550 ;
        RECT 18.270 16.490 18.630 16.990 ;
        RECT 18.335 14.550 18.565 16.490 ;
        RECT 18.870 14.390 19.310 18.710 ;
        RECT 19.625 15.610 19.855 18.550 ;
        RECT 19.550 14.610 19.930 15.610 ;
        RECT 19.625 14.550 19.855 14.610 ;
        RECT 20.150 14.390 20.590 18.710 ;
        RECT 20.915 18.490 21.145 18.550 ;
        RECT 20.820 17.490 21.240 18.490 ;
        RECT 20.915 14.550 21.145 17.490 ;
        RECT 21.455 14.390 21.895 18.710 ;
        RECT 22.415 18.695 23.435 18.710 ;
        RECT 22.205 15.610 22.435 18.550 ;
        RECT 22.130 14.610 22.510 15.610 ;
        RECT 22.205 14.550 22.435 14.610 ;
        RECT 22.730 14.390 23.170 18.695 ;
        RECT 23.495 16.985 23.725 18.550 ;
        RECT 23.430 16.485 23.790 16.985 ;
        RECT 23.495 14.550 23.725 16.485 ;
        RECT 24.005 14.390 24.535 18.710 ;
        RECT 25.280 18.695 26.015 18.710 ;
        RECT 24.785 15.610 25.015 18.550 ;
        RECT 24.720 14.610 25.080 15.610 ;
        RECT 24.785 14.550 25.015 14.610 ;
        RECT 25.280 14.390 25.810 18.695 ;
        RECT 26.075 16.985 26.305 18.550 ;
        RECT 26.010 16.485 26.370 16.985 ;
        RECT 26.075 14.550 26.305 16.485 ;
        RECT 26.630 14.390 27.070 18.710 ;
        RECT 27.365 15.610 27.595 18.550 ;
        RECT 27.290 14.610 27.670 15.610 ;
        RECT 27.365 14.550 27.595 14.610 ;
        RECT 27.910 14.390 28.350 18.710 ;
        RECT 28.655 18.490 28.885 18.550 ;
        RECT 28.560 17.490 28.980 18.490 ;
        RECT 28.655 14.550 28.885 17.490 ;
        RECT 29.205 14.390 29.645 18.710 ;
        RECT 30.155 18.695 31.175 18.710 ;
        RECT 31.770 18.695 32.465 18.710 ;
        RECT 29.945 15.610 30.175 18.550 ;
        RECT 29.870 14.610 30.250 15.610 ;
        RECT 29.945 14.550 30.175 14.610 ;
        RECT 30.505 14.390 30.945 18.695 ;
        RECT 31.235 16.985 31.465 18.550 ;
        RECT 31.170 16.485 31.530 16.985 ;
        RECT 31.235 14.550 31.465 16.485 ;
        RECT 31.770 14.390 32.210 18.695 ;
        RECT 32.525 15.610 32.755 18.550 ;
        RECT 32.460 14.610 32.820 15.610 ;
        RECT 32.525 14.550 32.755 14.610 ;
        RECT 1.845 14.160 2.805 14.390 ;
        RECT 3.135 14.160 7.965 14.390 ;
        RECT 8.295 14.160 10.545 14.390 ;
        RECT 10.875 14.160 15.705 14.390 ;
        RECT 16.035 14.160 18.285 14.390 ;
        RECT 18.615 14.160 23.445 14.390 ;
        RECT 23.775 14.160 26.025 14.390 ;
        RECT 26.355 14.160 31.185 14.390 ;
        RECT 31.515 14.160 32.475 14.390 ;
        RECT 1.385 12.725 33.215 13.345 ;
        RECT 1.350 12.000 4.105 12.540 ;
        RECT 5.885 11.615 6.485 11.675 ;
        RECT 0.920 10.150 5.140 10.410 ;
        RECT 0.650 9.450 1.310 9.510 ;
        RECT 0.630 7.055 1.330 9.450 ;
        RECT 2.090 7.360 5.140 10.150 ;
        RECT 0.650 6.995 1.310 7.055 ;
        RECT 1.105 5.795 5.350 6.595 ;
        RECT 5.865 6.400 6.505 11.615 ;
        RECT 10.360 8.625 37.515 9.640 ;
        RECT 11.275 8.030 17.395 8.260 ;
        RECT 17.725 8.030 23.845 8.260 ;
        RECT 24.175 8.030 30.295 8.260 ;
        RECT 30.625 8.030 36.745 8.260 ;
        RECT 10.995 7.810 11.225 7.870 ;
        RECT 10.930 7.510 11.290 7.810 ;
        RECT 10.995 6.870 11.225 7.510 ;
        RECT 11.580 6.710 11.915 8.030 ;
        RECT 12.285 7.810 12.515 7.870 ;
        RECT 12.220 7.510 12.580 7.810 ;
        RECT 12.285 6.870 12.515 7.510 ;
        RECT 12.870 6.710 13.205 8.030 ;
        RECT 13.575 7.230 13.805 8.030 ;
        RECT 13.510 6.710 13.870 7.230 ;
        RECT 14.180 6.710 14.515 8.030 ;
        RECT 14.865 7.810 15.095 7.870 ;
        RECT 14.800 7.510 15.160 7.810 ;
        RECT 14.865 6.870 15.095 7.510 ;
        RECT 15.465 6.710 15.800 8.030 ;
        RECT 16.155 7.230 16.385 8.030 ;
        RECT 16.090 6.710 16.450 7.230 ;
        RECT 16.765 6.710 17.100 8.030 ;
        RECT 17.445 7.810 17.675 7.870 ;
        RECT 17.380 7.510 17.740 7.810 ;
        RECT 17.445 6.870 17.675 7.510 ;
        RECT 18.025 6.710 18.360 8.030 ;
        RECT 18.735 7.810 18.965 7.870 ;
        RECT 18.670 7.510 19.030 7.810 ;
        RECT 18.735 6.870 18.965 7.510 ;
        RECT 19.295 6.710 19.630 8.030 ;
        RECT 20.025 7.230 20.255 8.030 ;
        RECT 19.960 6.710 20.320 7.230 ;
        RECT 20.600 6.710 20.935 8.030 ;
        RECT 21.315 7.810 21.545 7.870 ;
        RECT 21.250 7.510 21.610 7.810 ;
        RECT 21.315 6.870 21.545 7.510 ;
        RECT 21.865 6.710 22.200 8.030 ;
        RECT 22.605 7.230 22.835 8.030 ;
        RECT 22.540 6.710 22.900 7.230 ;
        RECT 23.175 6.710 23.510 8.030 ;
        RECT 23.895 7.810 24.125 7.870 ;
        RECT 23.830 7.510 24.190 7.810 ;
        RECT 23.895 6.870 24.125 7.510 ;
        RECT 24.465 6.710 24.800 8.030 ;
        RECT 25.185 7.810 25.415 7.870 ;
        RECT 25.120 7.510 25.480 7.810 ;
        RECT 25.185 6.870 25.415 7.510 ;
        RECT 25.750 6.710 26.085 8.030 ;
        RECT 26.475 7.230 26.705 8.030 ;
        RECT 26.410 6.710 26.770 7.230 ;
        RECT 27.055 6.710 27.390 8.030 ;
        RECT 27.765 7.810 27.995 7.870 ;
        RECT 27.700 7.510 28.060 7.810 ;
        RECT 27.765 6.870 27.995 7.510 ;
        RECT 28.350 6.710 28.685 8.030 ;
        RECT 29.055 7.230 29.285 8.030 ;
        RECT 28.990 6.710 29.350 7.230 ;
        RECT 29.600 6.710 29.935 8.030 ;
        RECT 30.345 7.810 30.575 7.870 ;
        RECT 30.280 7.510 30.640 7.810 ;
        RECT 30.345 6.870 30.575 7.510 ;
        RECT 30.900 6.710 31.235 8.030 ;
        RECT 31.635 7.810 31.865 7.870 ;
        RECT 31.570 7.510 31.930 7.810 ;
        RECT 31.635 6.870 31.865 7.510 ;
        RECT 32.210 6.710 32.545 8.030 ;
        RECT 32.925 7.230 33.155 8.030 ;
        RECT 32.860 6.710 33.220 7.230 ;
        RECT 33.510 6.710 33.845 8.030 ;
        RECT 34.215 7.810 34.445 7.870 ;
        RECT 34.150 7.510 34.510 7.810 ;
        RECT 34.215 6.870 34.445 7.510 ;
        RECT 34.805 6.710 35.140 8.030 ;
        RECT 35.505 7.230 35.735 8.030 ;
        RECT 35.440 6.710 35.800 7.230 ;
        RECT 36.140 6.710 36.475 8.030 ;
        RECT 36.795 7.810 37.025 7.870 ;
        RECT 36.730 7.510 37.090 7.810 ;
        RECT 36.795 7.230 37.025 7.510 ;
        RECT 36.730 6.930 37.090 7.230 ;
        RECT 36.795 6.870 37.025 6.930 ;
        RECT 11.275 6.480 17.395 6.710 ;
        RECT 17.725 6.480 23.845 6.710 ;
        RECT 24.175 6.480 30.295 6.710 ;
        RECT 30.625 6.480 36.745 6.710 ;
        RECT 5.885 6.340 6.485 6.400 ;
        RECT 1.300 4.365 3.195 4.470 ;
        RECT 3.570 4.365 5.465 4.470 ;
        RECT 8.765 4.365 37.095 4.370 ;
        RECT 0.975 4.140 37.095 4.365 ;
        RECT 0.975 4.135 12.005 4.140 ;
        RECT 0.975 3.430 1.205 4.135 ;
        RECT 1.550 3.225 2.960 4.135 ;
        RECT 3.265 3.870 3.495 3.930 ;
        RECT 3.200 3.490 3.560 3.870 ;
        RECT 3.265 3.430 3.495 3.490 ;
        RECT 3.785 3.225 5.195 4.135 ;
        RECT 5.555 3.430 5.785 4.135 ;
        RECT 6.600 3.870 6.830 3.930 ;
        RECT 1.255 2.995 3.215 3.225 ;
        RECT 3.545 2.995 5.505 3.225 ;
        RECT 6.505 3.170 6.925 3.870 ;
        RECT 6.600 2.930 6.830 3.170 ;
        RECT 7.095 2.725 7.685 4.135 ;
        RECT 7.890 3.690 8.120 3.930 ;
        RECT 7.825 2.990 8.185 3.690 ;
        RECT 7.890 2.930 8.120 2.990 ;
        RECT 8.355 2.725 8.945 4.135 ;
        RECT 9.180 3.870 9.410 3.930 ;
        RECT 9.085 3.170 9.505 3.870 ;
        RECT 12.575 3.610 12.805 3.935 ;
        RECT 9.180 2.930 9.410 3.170 ;
        RECT 12.510 2.995 12.870 3.610 ;
        RECT 12.575 2.935 12.805 2.995 ;
        RECT 13.105 2.730 14.500 4.140 ;
        RECT 14.865 3.875 15.095 3.935 ;
        RECT 14.800 3.310 15.160 3.875 ;
        RECT 19.025 3.610 19.255 3.935 ;
        RECT 14.865 2.935 15.095 3.310 ;
        RECT 18.960 2.995 19.320 3.610 ;
        RECT 19.025 2.935 19.255 2.995 ;
        RECT 19.595 2.730 20.990 4.140 ;
        RECT 21.315 3.875 21.545 3.935 ;
        RECT 21.250 3.310 21.610 3.875 ;
        RECT 25.475 3.610 25.705 3.935 ;
        RECT 21.315 2.935 21.545 3.310 ;
        RECT 25.410 2.995 25.770 3.610 ;
        RECT 25.475 2.935 25.705 2.995 ;
        RECT 26.000 2.730 27.395 4.140 ;
        RECT 27.765 3.875 27.995 3.935 ;
        RECT 27.700 3.310 28.060 3.875 ;
        RECT 31.925 3.615 32.155 3.935 ;
        RECT 27.765 2.935 27.995 3.310 ;
        RECT 31.860 2.995 32.220 3.615 ;
        RECT 31.925 2.935 32.155 2.995 ;
        RECT 32.550 2.730 33.945 4.140 ;
        RECT 34.215 3.875 34.445 3.935 ;
        RECT 34.150 3.260 34.510 3.875 ;
        RECT 34.830 3.610 35.060 3.935 ;
        RECT 34.215 2.935 34.445 3.260 ;
        RECT 34.765 2.995 35.125 3.610 ;
        RECT 34.830 2.935 35.060 2.995 ;
        RECT 35.430 2.730 36.825 4.140 ;
        RECT 37.120 3.875 37.350 3.935 ;
        RECT 37.055 3.260 37.415 3.875 ;
        RECT 37.120 2.935 37.350 3.260 ;
        RECT 6.880 2.495 7.840 2.725 ;
        RECT 8.170 2.495 9.130 2.725 ;
        RECT 12.855 2.500 14.815 2.730 ;
        RECT 19.305 2.500 21.265 2.730 ;
        RECT 25.755 2.500 27.715 2.730 ;
        RECT 32.205 2.500 34.165 2.730 ;
        RECT 35.110 2.500 37.070 2.730 ;
        RECT 5.025 2.225 10.075 2.235 ;
        RECT 0.060 1.505 10.075 2.225 ;
        RECT 30.970 1.670 31.260 1.690 ;
        RECT 5.025 1.500 10.075 1.505 ;
        RECT 0.065 0.370 10.080 1.170 ;
        RECT 12.510 0.915 37.655 1.670 ;
        RECT 30.970 0.895 31.260 0.915 ;
      LAYER met2 ;
        RECT -0.260 27.575 33.375 28.070 ;
        RECT -0.250 27.565 33.375 27.575 ;
        RECT -0.260 27.100 33.375 27.565 ;
        RECT 0.500 13.365 0.770 27.100 ;
        RECT 1.520 24.845 1.840 25.945 ;
        RECT 5.420 24.845 5.680 27.100 ;
        RECT 9.260 24.845 9.580 25.945 ;
        RECT 13.160 24.845 13.420 27.100 ;
        RECT 17.000 24.845 17.320 25.945 ;
        RECT 20.895 24.845 21.155 27.100 ;
        RECT 24.740 24.845 25.060 25.945 ;
        RECT 28.640 24.845 28.900 27.100 ;
        RECT 32.480 24.845 32.800 25.945 ;
        RECT 12.485 24.185 12.745 24.190 ;
        RECT 21.520 24.185 21.780 24.190 ;
        RECT 27.975 24.185 28.235 24.200 ;
        RECT 29.285 24.185 29.545 24.190 ;
        RECT 4.130 23.585 34.170 24.185 ;
        RECT 13.795 23.580 14.055 23.585 ;
        RECT 20.260 23.575 20.520 23.585 ;
        RECT 2.830 21.965 3.110 23.065 ;
        RECT 7.990 21.965 8.270 23.065 ;
        RECT 10.570 21.965 10.850 23.065 ;
        RECT 15.730 21.965 16.010 23.065 ;
        RECT 18.310 21.965 18.590 23.065 ;
        RECT 23.470 21.965 23.750 23.065 ;
        RECT 26.050 21.965 26.330 23.065 ;
        RECT 31.210 21.965 31.490 23.065 ;
        RECT 3.535 21.500 4.035 21.860 ;
        RECT 6.115 21.500 6.615 21.860 ;
        RECT 11.115 21.500 11.775 21.860 ;
        RECT 13.855 21.500 14.355 21.860 ;
        RECT 18.885 21.500 19.515 21.860 ;
        RECT 21.595 21.500 22.095 21.860 ;
        RECT 26.630 21.500 27.255 21.860 ;
        RECT 29.335 21.500 29.835 21.860 ;
        RECT 31.915 21.500 32.415 21.860 ;
        RECT 3.775 20.730 4.035 21.500 ;
        RECT 3.775 20.370 4.275 20.730 ;
        RECT 6.355 20.005 6.615 21.500 ;
        RECT 11.515 20.730 11.775 21.500 ;
        RECT 7.645 20.370 8.145 20.730 ;
        RECT 11.515 20.370 12.015 20.730 ;
        RECT 2.485 19.645 2.985 20.005 ;
        RECT 6.355 19.645 6.855 20.005 ;
        RECT 2.485 19.005 2.745 19.645 ;
        RECT 7.645 19.005 7.905 20.370 ;
        RECT 14.095 20.005 14.355 21.500 ;
        RECT 19.255 20.730 19.515 21.500 ;
        RECT 15.385 20.370 15.885 20.730 ;
        RECT 19.255 20.370 19.755 20.730 ;
        RECT 10.225 19.645 10.725 20.005 ;
        RECT 14.095 19.645 14.595 20.005 ;
        RECT 10.225 19.005 10.485 19.645 ;
        RECT 15.385 19.005 15.645 20.370 ;
        RECT 21.835 20.005 22.095 21.500 ;
        RECT 26.995 20.730 27.255 21.500 ;
        RECT 23.125 20.370 23.625 20.730 ;
        RECT 26.995 20.370 27.495 20.730 ;
        RECT 17.965 19.645 18.465 20.005 ;
        RECT 21.835 19.645 22.335 20.005 ;
        RECT 17.965 19.005 18.225 19.645 ;
        RECT 23.125 19.005 23.385 20.370 ;
        RECT 29.575 20.005 29.835 21.500 ;
        RECT 32.155 20.730 32.415 21.500 ;
        RECT 30.865 20.370 31.365 20.730 ;
        RECT 32.155 20.370 32.655 20.730 ;
        RECT 25.705 19.645 26.205 20.005 ;
        RECT 29.575 19.645 30.075 20.005 ;
        RECT 25.705 19.005 25.965 19.645 ;
        RECT 30.865 19.005 31.125 20.370 ;
        RECT 32.155 19.645 32.655 20.005 ;
        RECT 32.155 19.005 32.415 19.645 ;
        RECT 2.245 18.645 2.745 19.005 ;
        RECT 6.905 18.645 7.905 19.005 ;
        RECT 9.985 18.645 10.485 19.005 ;
        RECT 14.725 18.645 15.645 19.005 ;
        RECT 17.725 18.645 18.225 19.005 ;
        RECT 22.465 18.645 23.385 19.005 ;
        RECT 25.465 18.645 25.965 19.005 ;
        RECT 30.205 18.645 31.125 19.005 ;
        RECT 31.915 18.645 32.415 19.005 ;
        RECT 5.390 17.440 5.710 18.540 ;
        RECT 13.130 17.440 13.450 18.540 ;
        RECT 20.870 17.440 21.190 18.540 ;
        RECT 28.610 17.440 28.930 18.540 ;
        RECT 8.615 17.035 8.875 17.040 ;
        RECT 9.895 17.035 10.155 17.045 ;
        RECT 18.320 17.035 18.580 17.040 ;
        RECT 31.850 17.035 32.110 17.045 ;
        RECT 33.570 17.035 34.170 23.585 ;
        RECT 2.105 16.435 34.170 17.035 ;
        RECT 2.225 16.425 2.485 16.435 ;
        RECT 17.635 16.425 17.895 16.435 ;
        RECT 24.115 16.425 24.375 16.435 ;
        RECT 1.550 13.365 1.810 15.660 ;
        RECT 4.120 14.565 4.400 15.665 ;
        RECT 6.700 14.560 6.980 15.660 ;
        RECT 9.290 13.365 9.550 15.660 ;
        RECT 11.860 14.560 12.140 15.660 ;
        RECT 14.440 14.560 14.720 15.660 ;
        RECT 17.030 13.365 17.290 15.660 ;
        RECT 19.600 14.560 19.880 15.660 ;
        RECT 22.180 14.560 22.460 15.660 ;
        RECT 24.770 13.365 25.030 15.660 ;
        RECT 27.340 14.560 27.620 15.660 ;
        RECT 29.920 14.560 30.200 15.660 ;
        RECT 32.510 13.365 32.770 15.660 ;
        RECT 0.500 13.095 33.155 13.365 ;
        RECT 1.385 12.705 33.155 13.095 ;
        RECT 1.385 11.980 4.045 12.705 ;
        RECT 0.605 6.700 1.410 9.510 ;
        RECT 4.580 7.335 4.950 10.435 ;
        RECT 5.805 6.700 6.575 12.705 ;
        RECT 9.955 8.605 37.455 9.660 ;
        RECT 7.060 7.860 7.870 7.900 ;
        RECT 7.030 7.460 11.240 7.860 ;
        RECT 12.270 7.460 17.690 7.860 ;
        RECT 18.720 7.460 24.140 7.860 ;
        RECT 25.170 7.460 30.590 7.860 ;
        RECT 31.620 7.460 37.040 7.860 ;
        RECT 7.060 7.430 7.870 7.460 ;
        RECT 13.560 6.880 16.400 7.280 ;
        RECT 20.010 6.880 22.850 7.280 ;
        RECT 26.460 6.880 29.300 7.280 ;
        RECT 32.910 6.880 35.750 7.280 ;
        RECT 0.605 5.750 6.575 6.700 ;
        RECT 1.350 4.095 3.145 4.520 ;
        RECT 3.620 4.095 5.415 4.520 ;
        RECT 1.950 2.245 2.210 2.340 ;
        RECT 3.250 2.245 3.510 3.920 ;
        RECT 6.555 3.120 6.875 3.920 ;
        RECT 7.875 2.255 8.135 3.740 ;
        RECT 9.135 3.120 9.455 3.920 ;
        RECT 5.085 2.245 10.015 2.255 ;
        RECT 0.120 1.915 10.015 2.245 ;
        RECT 0.115 1.515 10.015 1.915 ;
        RECT 12.560 1.690 12.820 3.660 ;
        RECT 14.850 3.260 15.110 6.880 ;
        RECT 19.010 1.690 19.270 3.660 ;
        RECT 21.300 3.260 21.560 6.880 ;
        RECT 25.460 1.690 25.720 3.660 ;
        RECT 27.750 3.260 28.010 6.880 ;
        RECT 31.910 1.720 32.170 3.665 ;
        RECT 34.200 3.215 34.460 6.880 ;
        RECT 36.780 5.315 37.040 7.460 ;
        RECT 36.780 5.195 38.335 5.315 ;
        RECT 36.780 5.185 38.325 5.195 ;
        RECT 36.780 5.070 38.335 5.185 ;
        RECT 34.815 1.720 35.075 3.660 ;
        RECT 37.105 3.210 37.365 5.070 ;
        RECT 38.150 5.055 38.335 5.070 ;
        RECT 30.835 1.690 38.565 1.720 ;
        RECT 11.705 1.515 38.565 1.690 ;
        RECT 0.115 1.195 38.565 1.515 ;
        RECT -0.110 1.170 38.565 1.195 ;
        RECT -0.165 0.970 38.565 1.170 ;
        RECT -0.165 0.960 38.550 0.970 ;
        RECT 38.560 0.960 38.565 0.970 ;
        RECT -0.165 0.350 38.565 0.960 ;
        RECT -0.110 0.180 38.565 0.350 ;
      LAYER met3 ;
        RECT 1.470 24.870 1.890 25.920 ;
        RECT 9.210 24.870 9.630 25.920 ;
        RECT 16.950 24.870 17.370 25.920 ;
        RECT 24.690 24.870 25.110 25.920 ;
        RECT 32.430 24.870 32.850 25.920 ;
        RECT 2.780 22.370 3.160 23.040 ;
        RECT 7.940 22.370 8.320 23.040 ;
        RECT 10.520 22.370 10.900 23.040 ;
        RECT 15.680 22.370 16.060 23.040 ;
        RECT 18.260 22.370 18.640 23.040 ;
        RECT 23.420 22.370 23.800 23.040 ;
        RECT 26.000 22.370 26.380 23.040 ;
        RECT 31.160 22.370 31.540 23.040 ;
        RECT 0.830 22.000 31.540 22.370 ;
        RECT 0.830 14.965 1.200 22.000 ;
        RECT 2.780 21.990 3.160 22.000 ;
        RECT 7.940 21.990 8.320 22.000 ;
        RECT 10.520 21.990 10.900 22.000 ;
        RECT 15.680 21.990 16.060 22.000 ;
        RECT 18.260 21.990 18.640 22.000 ;
        RECT 23.420 21.990 23.800 22.000 ;
        RECT 26.000 21.990 26.380 22.000 ;
        RECT 30.840 21.990 31.540 22.000 ;
        RECT 5.340 17.465 5.760 18.515 ;
        RECT 13.080 17.465 13.500 18.515 ;
        RECT 20.820 17.465 21.240 18.515 ;
        RECT 28.560 17.465 28.980 18.515 ;
        RECT 4.070 14.965 4.450 15.640 ;
        RECT 6.650 14.965 7.030 15.635 ;
        RECT 11.810 14.965 12.190 15.635 ;
        RECT 14.390 14.965 14.770 15.635 ;
        RECT 19.550 14.965 19.930 15.635 ;
        RECT 22.130 14.965 22.510 15.635 ;
        RECT 27.290 14.965 27.670 15.635 ;
        RECT 29.870 14.965 30.250 15.635 ;
        RECT 0.830 14.585 30.250 14.965 ;
        RECT 4.530 7.360 5.000 10.410 ;
        RECT 7.030 7.875 7.410 14.585 ;
        RECT 7.010 7.455 7.920 7.875 ;
        RECT 1.300 4.120 3.195 4.495 ;
        RECT 3.570 4.120 5.465 4.495 ;
        RECT 6.505 3.145 6.925 3.895 ;
        RECT 9.085 3.145 9.505 3.895 ;
      LAYER met4 ;
        RECT 0.100 25.520 32.805 25.900 ;
        RECT 0.100 22.245 0.480 25.520 ;
        RECT 1.515 24.890 1.845 25.520 ;
        RECT 9.255 24.890 9.585 25.520 ;
        RECT 16.995 24.890 17.325 25.520 ;
        RECT 24.735 24.890 25.065 25.520 ;
        RECT 32.475 24.890 32.805 25.520 ;
        RECT -0.840 21.860 0.480 22.245 ;
        RECT -0.840 4.495 -0.460 21.860 ;
        RECT 0.100 18.495 0.480 21.860 ;
        RECT 0.100 18.115 28.935 18.495 ;
        RECT 5.385 17.485 5.715 18.115 ;
        RECT 13.125 17.485 13.455 18.115 ;
        RECT 20.865 17.485 21.195 18.115 ;
        RECT 28.605 17.485 28.935 18.115 ;
        RECT 4.575 7.740 4.955 10.390 ;
        RECT 4.575 7.360 8.185 7.740 ;
        RECT 7.855 5.400 8.185 7.360 ;
        RECT 6.550 5.020 9.460 5.400 ;
        RECT -0.840 4.130 5.605 4.495 ;
        RECT 6.550 3.165 6.880 5.020 ;
        RECT 9.130 3.165 9.460 5.020 ;
  END
END BGR_BJT_final
END LIBRARY

