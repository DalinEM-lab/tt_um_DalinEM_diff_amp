magic
tech sky130A
magscale 1 2
timestamp 1741231714
<< nwell >>
rect -10291 3942 -2281 5417
rect -1833 -136 780 7623
rect 3203 -7 5209 1831
rect 7129 83 12023 2517
rect 11629 -1147 12447 -189
rect 3054 -4162 3689 -2789
rect 3038 -5458 3676 -4666
rect 3038 -6748 3676 -5956
rect 3038 -8038 3676 -7246
rect 3045 -9163 3677 -8332
rect 3044 -10343 3677 -9163
rect 3044 -10347 3676 -10343
<< pwell >>
rect -10287 428 -9267 1820
rect -9027 -103 -3500 3452
rect -8943 -137 -8920 -103
rect -8826 -137 -3593 -135
rect 8505 -2337 10641 -52
rect -1564 -8169 1550 -3519
rect -1564 -8201 -320 -8169
rect -316 -8170 1550 -8169
rect -316 -8201 -270 -8170
rect -1564 -8203 -270 -8201
rect -267 -8203 1550 -8170
rect -1564 -10361 1550 -8203
rect 2146 -8449 2993 -2775
rect 8830 -3535 10350 -2485
rect 11109 -2605 12513 -2203
rect 1596 -9120 2936 -8967
rect 1596 -10154 1749 -9120
rect 2783 -10154 2936 -9120
rect 1596 -10307 2936 -10154
<< nbase >>
rect 1749 -10154 2783 -9120
<< nmos >>
rect -10077 624 -9477 1624
rect 9040 -2981 10140 -2681
rect 9040 -3339 10140 -3039
<< pmos >>
rect 3399 212 3759 1612
rect 3817 212 4177 1612
rect 4235 212 4595 1612
rect 4653 212 5013 1612
<< pmoslvt >>
rect -9902 4707 -6302 5067
rect -6244 4707 -2644 5067
rect -9902 4219 -6302 4579
rect -6244 4219 -2644 4579
rect -1430 4143 -1050 7143
rect -992 4143 -612 7143
rect -554 4143 -174 7143
rect -116 4143 264 7143
rect -1430 166 -1050 3166
rect -992 166 -612 3166
rect -554 166 -174 3166
rect -116 166 264 3166
rect 7492 1657 8492 2157
rect 8550 1657 9550 2157
rect 9608 1657 10608 2157
rect 10666 1657 11666 2157
rect 7492 495 8492 995
rect 8550 495 9550 995
rect 9608 495 10608 995
rect 10666 495 11666 995
rect 11825 -928 11895 -408
rect 12181 -928 12251 -408
rect 3257 -3391 3457 -2991
rect 3257 -3972 3457 -3572
rect 3257 -5262 3457 -4862
rect 3257 -6552 3457 -6152
rect 3257 -7842 3457 -7442
rect 3257 -8730 3457 -8530
rect 3257 -8988 3457 -8788
rect 3257 -9655 3357 -9255
rect 3257 -10113 3357 -9713
<< nmoslvt >>
rect -8692 1995 -6292 3195
rect -6234 1995 -3834 3195
rect -8693 120 -6293 1320
rect -6235 120 -3835 1320
rect -1420 -1160 460 -860
rect 518 -1160 2398 -860
rect 2456 -1160 4336 -860
rect 4394 -1160 6274 -860
rect -1420 -1570 460 -1270
rect 518 -1570 2398 -1270
rect 2456 -1570 4336 -1270
rect 4394 -1570 6274 -1270
rect 8677 -890 9077 -290
rect 9135 -890 9535 -290
rect 9593 -890 9993 -290
rect 10051 -890 10451 -290
rect 8677 -2097 9077 -1497
rect 9135 -2097 9535 -1497
rect 9593 -2097 9993 -1497
rect 10051 -2097 10451 -1497
rect 11865 -1613 11895 -1413
rect 12221 -1613 12251 -1413
rect -1148 -4061 -348 -3861
rect 333 -4061 1133 -3861
rect -1148 -4319 -348 -4119
rect 333 -4319 1133 -4119
rect -1148 -4577 -348 -4377
rect 333 -4577 1133 -4377
rect -1148 -4835 -348 -4635
rect 333 -4835 1133 -4635
rect -1148 -5093 -348 -4893
rect 333 -5093 1133 -4893
rect -1148 -5351 -348 -5151
rect 333 -5351 1133 -5151
rect -1148 -5609 -348 -5409
rect 333 -5609 1133 -5409
rect -1148 -5867 -348 -5667
rect 333 -5867 1133 -5667
rect -1148 -6125 -348 -5925
rect 333 -6125 1133 -5925
rect -1148 -6383 -348 -6183
rect 333 -6383 1133 -6183
rect -1148 -6641 -348 -6441
rect 333 -6641 1133 -6441
rect -1148 -6899 -348 -6699
rect 333 -6899 1133 -6699
rect -1148 -7157 -348 -6957
rect 333 -7157 1133 -6957
rect -1148 -7415 -348 -7215
rect 333 -7415 1133 -7215
rect -1148 -7673 -348 -7473
rect 333 -7673 1133 -7473
rect -1148 -7931 -348 -7731
rect 333 -7931 1133 -7731
rect -1148 -8189 -348 -7989
rect 333 -8189 1133 -7989
rect -1148 -8447 -348 -8247
rect 333 -8447 1133 -8247
rect -1148 -8705 -348 -8505
rect 333 -8705 1133 -8505
rect -1148 -8963 -348 -8763
rect 333 -8963 1133 -8763
rect -1148 -9221 -348 -9021
rect 333 -9221 1133 -9021
rect -1148 -9479 -348 -9279
rect 333 -9479 1133 -9279
rect -1148 -9737 -348 -9537
rect 333 -9737 1133 -9537
rect -1148 -9995 -348 -9795
rect 333 -9995 1133 -9795
rect 2470 -3256 2670 -3056
rect 2470 -3514 2670 -3314
rect 2470 -3772 2670 -3572
rect 2470 -4030 2670 -3830
rect 2470 -4288 2670 -4088
rect 2470 -4546 2670 -4346
rect 2470 -4804 2670 -4604
rect 2470 -5062 2670 -4862
rect 2470 -5320 2670 -5120
rect 2470 -5578 2670 -5378
rect 2470 -5836 2670 -5636
rect 2470 -6094 2670 -5894
rect 2470 -6352 2670 -6152
rect 2470 -6610 2670 -6410
rect 2470 -6868 2670 -6668
rect 2470 -7126 2670 -6926
rect 2470 -7384 2670 -7184
rect 2470 -7642 2670 -7442
rect 2470 -7900 2670 -7700
rect 2470 -8158 2670 -7958
<< ndiff >>
rect -10077 1670 -9477 1682
rect -10077 1636 -10065 1670
rect -9489 1636 -9477 1670
rect -10077 1624 -9477 1636
rect -10077 612 -9477 624
rect -10077 578 -10065 612
rect -9489 578 -9477 612
rect -10077 566 -9477 578
rect -8750 3183 -8692 3195
rect -8750 2007 -8738 3183
rect -8704 2007 -8692 3183
rect -8750 1995 -8692 2007
rect -6292 3183 -6234 3195
rect -6292 2007 -6280 3183
rect -6246 2007 -6234 3183
rect -6292 1995 -6234 2007
rect -3834 3183 -3776 3195
rect -3834 2007 -3822 3183
rect -3788 2007 -3776 3183
rect -3834 1995 -3776 2007
rect -8751 1308 -8693 1320
rect -8751 132 -8739 1308
rect -8705 132 -8693 1308
rect -8751 120 -8693 132
rect -6293 1308 -6235 1320
rect -6293 132 -6281 1308
rect -6247 132 -6235 1308
rect -6293 120 -6235 132
rect -3835 1308 -3777 1320
rect -3835 132 -3823 1308
rect -3789 132 -3777 1308
rect -3835 120 -3777 132
rect -1478 -872 -1420 -860
rect -1478 -1148 -1466 -872
rect -1432 -1148 -1420 -872
rect -1478 -1160 -1420 -1148
rect 460 -872 518 -860
rect 460 -1148 472 -872
rect 506 -1148 518 -872
rect 460 -1160 518 -1148
rect 2398 -872 2456 -860
rect 2398 -1148 2410 -872
rect 2444 -1148 2456 -872
rect 2398 -1160 2456 -1148
rect 4336 -872 4394 -860
rect 4336 -1148 4348 -872
rect 4382 -1148 4394 -872
rect 4336 -1160 4394 -1148
rect 6274 -872 6332 -860
rect 6274 -1148 6286 -872
rect 6320 -1148 6332 -872
rect 6274 -1160 6332 -1148
rect -1478 -1282 -1420 -1270
rect -1478 -1558 -1466 -1282
rect -1432 -1558 -1420 -1282
rect -1478 -1570 -1420 -1558
rect 460 -1282 518 -1270
rect 460 -1558 472 -1282
rect 506 -1558 518 -1282
rect 460 -1570 518 -1558
rect 2398 -1282 2456 -1270
rect 2398 -1558 2410 -1282
rect 2444 -1558 2456 -1282
rect 2398 -1570 2456 -1558
rect 4336 -1282 4394 -1270
rect 4336 -1558 4348 -1282
rect 4382 -1558 4394 -1282
rect 4336 -1570 4394 -1558
rect 6274 -1282 6332 -1270
rect 6274 -1558 6286 -1282
rect 6320 -1558 6332 -1282
rect 6274 -1570 6332 -1558
rect 8619 -302 8677 -290
rect 8619 -878 8631 -302
rect 8665 -878 8677 -302
rect 8619 -890 8677 -878
rect 9077 -302 9135 -290
rect 9077 -878 9089 -302
rect 9123 -878 9135 -302
rect 9077 -890 9135 -878
rect 9535 -302 9593 -290
rect 9535 -878 9547 -302
rect 9581 -878 9593 -302
rect 9535 -890 9593 -878
rect 9993 -302 10051 -290
rect 9993 -878 10005 -302
rect 10039 -878 10051 -302
rect 9993 -890 10051 -878
rect 10451 -302 10509 -290
rect 10451 -878 10463 -302
rect 10497 -878 10509 -302
rect 10451 -890 10509 -878
rect 8619 -1509 8677 -1497
rect 8619 -2085 8631 -1509
rect 8665 -2085 8677 -1509
rect 8619 -2097 8677 -2085
rect 9077 -1509 9135 -1497
rect 9077 -2085 9089 -1509
rect 9123 -2085 9135 -1509
rect 9077 -2097 9135 -2085
rect 9535 -1509 9593 -1497
rect 9535 -2085 9547 -1509
rect 9581 -2085 9593 -1509
rect 9535 -2097 9593 -2085
rect 9993 -1509 10051 -1497
rect 9993 -2085 10005 -1509
rect 10039 -2085 10051 -1509
rect 9993 -2097 10051 -2085
rect 10451 -1509 10509 -1497
rect 10451 -2085 10463 -1509
rect 10497 -2085 10509 -1509
rect 10451 -2097 10509 -2085
rect 11807 -1425 11865 -1413
rect 11807 -1601 11819 -1425
rect 11853 -1601 11865 -1425
rect 11807 -1613 11865 -1601
rect 11895 -1425 11953 -1413
rect 11895 -1601 11907 -1425
rect 11941 -1601 11953 -1425
rect 11895 -1613 11953 -1601
rect 12163 -1425 12221 -1413
rect 12163 -1601 12175 -1425
rect 12209 -1601 12221 -1425
rect 12163 -1613 12221 -1601
rect 12251 -1425 12309 -1413
rect 12251 -1601 12263 -1425
rect 12297 -1601 12309 -1425
rect 12251 -1613 12309 -1601
rect -1148 -3815 -348 -3803
rect -1148 -3849 -1136 -3815
rect -360 -3849 -348 -3815
rect -1148 -3861 -348 -3849
rect 333 -3815 1133 -3803
rect 333 -3849 345 -3815
rect 1121 -3849 1133 -3815
rect 333 -3861 1133 -3849
rect -1148 -4073 -348 -4061
rect -1148 -4107 -1136 -4073
rect -360 -4107 -348 -4073
rect -1148 -4119 -348 -4107
rect 333 -4073 1133 -4061
rect 333 -4107 345 -4073
rect 1121 -4107 1133 -4073
rect 333 -4119 1133 -4107
rect -1148 -4331 -348 -4319
rect -1148 -4365 -1136 -4331
rect -360 -4365 -348 -4331
rect -1148 -4377 -348 -4365
rect 333 -4331 1133 -4319
rect 333 -4365 345 -4331
rect 1121 -4365 1133 -4331
rect 333 -4377 1133 -4365
rect -1148 -4589 -348 -4577
rect -1148 -4623 -1136 -4589
rect -360 -4623 -348 -4589
rect -1148 -4635 -348 -4623
rect 333 -4589 1133 -4577
rect 333 -4623 345 -4589
rect 1121 -4623 1133 -4589
rect 333 -4635 1133 -4623
rect -1148 -4847 -348 -4835
rect -1148 -4881 -1136 -4847
rect -360 -4881 -348 -4847
rect -1148 -4893 -348 -4881
rect 333 -4847 1133 -4835
rect 333 -4881 345 -4847
rect 1121 -4881 1133 -4847
rect 333 -4893 1133 -4881
rect -1148 -5105 -348 -5093
rect -1148 -5139 -1136 -5105
rect -360 -5139 -348 -5105
rect -1148 -5151 -348 -5139
rect 333 -5105 1133 -5093
rect 333 -5139 345 -5105
rect 1121 -5139 1133 -5105
rect 333 -5151 1133 -5139
rect -1148 -5363 -348 -5351
rect -1148 -5397 -1136 -5363
rect -360 -5397 -348 -5363
rect -1148 -5409 -348 -5397
rect 333 -5363 1133 -5351
rect 333 -5397 345 -5363
rect 1121 -5397 1133 -5363
rect 333 -5409 1133 -5397
rect -1148 -5621 -348 -5609
rect -1148 -5655 -1136 -5621
rect -360 -5655 -348 -5621
rect -1148 -5667 -348 -5655
rect 333 -5621 1133 -5609
rect 333 -5655 345 -5621
rect 1121 -5655 1133 -5621
rect 333 -5667 1133 -5655
rect -1148 -5879 -348 -5867
rect -1148 -5913 -1136 -5879
rect -360 -5913 -348 -5879
rect -1148 -5925 -348 -5913
rect 333 -5879 1133 -5867
rect 333 -5913 345 -5879
rect 1121 -5913 1133 -5879
rect 333 -5925 1133 -5913
rect -1148 -6137 -348 -6125
rect -1148 -6171 -1136 -6137
rect -360 -6171 -348 -6137
rect -1148 -6183 -348 -6171
rect 333 -6137 1133 -6125
rect 333 -6171 345 -6137
rect 1121 -6171 1133 -6137
rect 333 -6183 1133 -6171
rect -1148 -6395 -348 -6383
rect -1148 -6429 -1136 -6395
rect -360 -6429 -348 -6395
rect -1148 -6441 -348 -6429
rect 333 -6395 1133 -6383
rect 333 -6429 345 -6395
rect 1121 -6429 1133 -6395
rect 333 -6441 1133 -6429
rect -1148 -6653 -348 -6641
rect -1148 -6687 -1136 -6653
rect -360 -6687 -348 -6653
rect -1148 -6699 -348 -6687
rect 333 -6653 1133 -6641
rect 333 -6687 345 -6653
rect 1121 -6687 1133 -6653
rect 333 -6699 1133 -6687
rect -1148 -6911 -348 -6899
rect -1148 -6945 -1136 -6911
rect -360 -6945 -348 -6911
rect -1148 -6957 -348 -6945
rect 333 -6911 1133 -6899
rect 333 -6945 345 -6911
rect 1121 -6945 1133 -6911
rect 333 -6957 1133 -6945
rect -1148 -7169 -348 -7157
rect -1148 -7203 -1136 -7169
rect -360 -7203 -348 -7169
rect -1148 -7215 -348 -7203
rect 333 -7169 1133 -7157
rect 333 -7203 345 -7169
rect 1121 -7203 1133 -7169
rect 333 -7215 1133 -7203
rect -1148 -7427 -348 -7415
rect -1148 -7461 -1136 -7427
rect -360 -7461 -348 -7427
rect -1148 -7473 -348 -7461
rect 333 -7427 1133 -7415
rect 333 -7461 345 -7427
rect 1121 -7461 1133 -7427
rect 333 -7473 1133 -7461
rect -1148 -7685 -348 -7673
rect -1148 -7719 -1136 -7685
rect -360 -7719 -348 -7685
rect -1148 -7731 -348 -7719
rect 333 -7685 1133 -7673
rect 333 -7719 345 -7685
rect 1121 -7719 1133 -7685
rect 333 -7731 1133 -7719
rect -1148 -7943 -348 -7931
rect -1148 -7977 -1136 -7943
rect -360 -7977 -348 -7943
rect -1148 -7989 -348 -7977
rect 333 -7943 1133 -7931
rect 333 -7977 345 -7943
rect 1121 -7977 1133 -7943
rect 333 -7989 1133 -7977
rect -1148 -8201 -348 -8189
rect -1148 -8235 -1136 -8201
rect -360 -8235 -348 -8201
rect -1148 -8247 -348 -8235
rect 333 -8201 1133 -8189
rect 333 -8235 345 -8201
rect 1121 -8235 1133 -8201
rect 333 -8247 1133 -8235
rect -1148 -8459 -348 -8447
rect -1148 -8493 -1136 -8459
rect -360 -8493 -348 -8459
rect -1148 -8505 -348 -8493
rect 333 -8459 1133 -8447
rect 333 -8493 345 -8459
rect 1121 -8493 1133 -8459
rect 333 -8505 1133 -8493
rect -1148 -8717 -348 -8705
rect -1148 -8751 -1136 -8717
rect -360 -8751 -348 -8717
rect -1148 -8763 -348 -8751
rect 333 -8717 1133 -8705
rect 333 -8751 345 -8717
rect 1121 -8751 1133 -8717
rect 333 -8763 1133 -8751
rect -1148 -8975 -348 -8963
rect -1148 -9009 -1136 -8975
rect -360 -9009 -348 -8975
rect -1148 -9021 -348 -9009
rect 333 -8975 1133 -8963
rect 333 -9009 345 -8975
rect 1121 -9009 1133 -8975
rect 333 -9021 1133 -9009
rect -1148 -9233 -348 -9221
rect -1148 -9267 -1136 -9233
rect -360 -9267 -348 -9233
rect -1148 -9279 -348 -9267
rect 333 -9233 1133 -9221
rect 333 -9267 345 -9233
rect 1121 -9267 1133 -9233
rect 333 -9279 1133 -9267
rect -1148 -9491 -348 -9479
rect -1148 -9525 -1136 -9491
rect -360 -9525 -348 -9491
rect -1148 -9537 -348 -9525
rect 333 -9491 1133 -9479
rect 333 -9525 345 -9491
rect 1121 -9525 1133 -9491
rect 333 -9537 1133 -9525
rect -1148 -9749 -348 -9737
rect -1148 -9783 -1136 -9749
rect -360 -9783 -348 -9749
rect -1148 -9795 -348 -9783
rect 333 -9749 1133 -9737
rect 333 -9783 345 -9749
rect 1121 -9783 1133 -9749
rect 333 -9795 1133 -9783
rect -1148 -10007 -348 -9995
rect -1148 -10041 -1136 -10007
rect -360 -10041 -348 -10007
rect -1148 -10053 -348 -10041
rect 333 -10007 1133 -9995
rect 333 -10041 345 -10007
rect 1121 -10041 1133 -10007
rect 333 -10053 1133 -10041
rect 2470 -3010 2670 -2998
rect 2470 -3044 2482 -3010
rect 2658 -3044 2670 -3010
rect 2470 -3056 2670 -3044
rect 2470 -3268 2670 -3256
rect 2470 -3302 2482 -3268
rect 2658 -3302 2670 -3268
rect 2470 -3314 2670 -3302
rect 2470 -3526 2670 -3514
rect 2470 -3560 2482 -3526
rect 2658 -3560 2670 -3526
rect 2470 -3572 2670 -3560
rect 2470 -3784 2670 -3772
rect 2470 -3818 2482 -3784
rect 2658 -3818 2670 -3784
rect 2470 -3830 2670 -3818
rect 2470 -4042 2670 -4030
rect 2470 -4076 2482 -4042
rect 2658 -4076 2670 -4042
rect 2470 -4088 2670 -4076
rect 2470 -4300 2670 -4288
rect 2470 -4334 2482 -4300
rect 2658 -4334 2670 -4300
rect 2470 -4346 2670 -4334
rect 2470 -4558 2670 -4546
rect 2470 -4592 2482 -4558
rect 2658 -4592 2670 -4558
rect 2470 -4604 2670 -4592
rect 2470 -4816 2670 -4804
rect 2470 -4850 2482 -4816
rect 2658 -4850 2670 -4816
rect 2470 -4862 2670 -4850
rect 2470 -5074 2670 -5062
rect 2470 -5108 2482 -5074
rect 2658 -5108 2670 -5074
rect 2470 -5120 2670 -5108
rect 2470 -5332 2670 -5320
rect 2470 -5366 2482 -5332
rect 2658 -5366 2670 -5332
rect 2470 -5378 2670 -5366
rect 2470 -5590 2670 -5578
rect 2470 -5624 2482 -5590
rect 2658 -5624 2670 -5590
rect 2470 -5636 2670 -5624
rect 2470 -5848 2670 -5836
rect 2470 -5882 2482 -5848
rect 2658 -5882 2670 -5848
rect 2470 -5894 2670 -5882
rect 2470 -6106 2670 -6094
rect 2470 -6140 2482 -6106
rect 2658 -6140 2670 -6106
rect 2470 -6152 2670 -6140
rect 2470 -6364 2670 -6352
rect 2470 -6398 2482 -6364
rect 2658 -6398 2670 -6364
rect 2470 -6410 2670 -6398
rect 2470 -6622 2670 -6610
rect 2470 -6656 2482 -6622
rect 2658 -6656 2670 -6622
rect 2470 -6668 2670 -6656
rect 2470 -6880 2670 -6868
rect 2470 -6914 2482 -6880
rect 2658 -6914 2670 -6880
rect 2470 -6926 2670 -6914
rect 2470 -7138 2670 -7126
rect 2470 -7172 2482 -7138
rect 2658 -7172 2670 -7138
rect 2470 -7184 2670 -7172
rect 2470 -7396 2670 -7384
rect 2470 -7430 2482 -7396
rect 2658 -7430 2670 -7396
rect 2470 -7442 2670 -7430
rect 2470 -7654 2670 -7642
rect 2470 -7688 2482 -7654
rect 2658 -7688 2670 -7654
rect 2470 -7700 2670 -7688
rect 2470 -7912 2670 -7900
rect 2470 -7946 2482 -7912
rect 2658 -7946 2670 -7912
rect 2470 -7958 2670 -7946
rect 2470 -8170 2670 -8158
rect 2470 -8204 2482 -8170
rect 2658 -8204 2670 -8170
rect 2470 -8216 2670 -8204
rect 9040 -2635 10140 -2623
rect 9040 -2669 9052 -2635
rect 10128 -2669 10140 -2635
rect 9040 -2681 10140 -2669
rect 9040 -2993 10140 -2981
rect 9040 -3027 9052 -2993
rect 10128 -3027 10140 -2993
rect 9040 -3039 10140 -3027
rect 9040 -3351 10140 -3339
rect 9040 -3385 9052 -3351
rect 10128 -3385 10140 -3351
rect 9040 -3397 10140 -3385
<< pdiff >>
rect -9960 5055 -9902 5067
rect -9960 4719 -9948 5055
rect -9914 4719 -9902 5055
rect -9960 4707 -9902 4719
rect -6302 5055 -6244 5067
rect -6302 4719 -6290 5055
rect -6256 4719 -6244 5055
rect -6302 4707 -6244 4719
rect -2644 5055 -2586 5067
rect -2644 4719 -2632 5055
rect -2598 4719 -2586 5055
rect -2644 4707 -2586 4719
rect -9960 4567 -9902 4579
rect -9960 4231 -9948 4567
rect -9914 4231 -9902 4567
rect -9960 4219 -9902 4231
rect -6302 4567 -6244 4579
rect -6302 4231 -6290 4567
rect -6256 4231 -6244 4567
rect -6302 4219 -6244 4231
rect -2644 4567 -2586 4579
rect -2644 4231 -2632 4567
rect -2598 4231 -2586 4567
rect -2644 4219 -2586 4231
rect -1488 7131 -1430 7143
rect -1488 4155 -1476 7131
rect -1442 4155 -1430 7131
rect -1488 4143 -1430 4155
rect -1050 7131 -992 7143
rect -1050 4155 -1038 7131
rect -1004 4155 -992 7131
rect -1050 4143 -992 4155
rect -612 7131 -554 7143
rect -612 4155 -600 7131
rect -566 4155 -554 7131
rect -612 4143 -554 4155
rect -174 7131 -116 7143
rect -174 4155 -162 7131
rect -128 4155 -116 7131
rect -174 4143 -116 4155
rect 264 7131 322 7143
rect 264 4155 276 7131
rect 310 4155 322 7131
rect 264 4143 322 4155
rect -1488 3154 -1430 3166
rect -1488 178 -1476 3154
rect -1442 178 -1430 3154
rect -1488 166 -1430 178
rect -1050 3154 -992 3166
rect -1050 178 -1038 3154
rect -1004 178 -992 3154
rect -1050 166 -992 178
rect -612 3154 -554 3166
rect -612 178 -600 3154
rect -566 178 -554 3154
rect -612 166 -554 178
rect -174 3154 -116 3166
rect -174 178 -162 3154
rect -128 178 -116 3154
rect -174 166 -116 178
rect 264 3154 322 3166
rect 264 178 276 3154
rect 310 178 322 3154
rect 264 166 322 178
rect 3341 1600 3399 1612
rect 3341 224 3353 1600
rect 3387 224 3399 1600
rect 3341 212 3399 224
rect 3759 1600 3817 1612
rect 3759 224 3771 1600
rect 3805 224 3817 1600
rect 3759 212 3817 224
rect 4177 1600 4235 1612
rect 4177 224 4189 1600
rect 4223 224 4235 1600
rect 4177 212 4235 224
rect 4595 1600 4653 1612
rect 4595 224 4607 1600
rect 4641 224 4653 1600
rect 4595 212 4653 224
rect 5013 1600 5071 1612
rect 5013 224 5025 1600
rect 5059 224 5071 1600
rect 5013 212 5071 224
rect 7434 2145 7492 2157
rect 7434 1669 7446 2145
rect 7480 1669 7492 2145
rect 7434 1657 7492 1669
rect 8492 2145 8550 2157
rect 8492 1669 8504 2145
rect 8538 1669 8550 2145
rect 8492 1657 8550 1669
rect 9550 2145 9608 2157
rect 9550 1669 9562 2145
rect 9596 1669 9608 2145
rect 9550 1657 9608 1669
rect 10608 2145 10666 2157
rect 10608 1669 10620 2145
rect 10654 1669 10666 2145
rect 10608 1657 10666 1669
rect 11666 2145 11724 2157
rect 11666 1669 11678 2145
rect 11712 1669 11724 2145
rect 11666 1657 11724 1669
rect 7434 983 7492 995
rect 7434 507 7446 983
rect 7480 507 7492 983
rect 7434 495 7492 507
rect 8492 983 8550 995
rect 8492 507 8504 983
rect 8538 507 8550 983
rect 8492 495 8550 507
rect 9550 983 9608 995
rect 9550 507 9562 983
rect 9596 507 9608 983
rect 9550 495 9608 507
rect 10608 983 10666 995
rect 10608 507 10620 983
rect 10654 507 10666 983
rect 10608 495 10666 507
rect 11666 983 11724 995
rect 11666 507 11678 983
rect 11712 507 11724 983
rect 11666 495 11724 507
rect 11767 -420 11825 -408
rect 11767 -916 11779 -420
rect 11813 -916 11825 -420
rect 11767 -928 11825 -916
rect 11895 -420 11953 -408
rect 11895 -916 11907 -420
rect 11941 -916 11953 -420
rect 11895 -928 11953 -916
rect 12123 -420 12181 -408
rect 12123 -916 12135 -420
rect 12169 -916 12181 -420
rect 12123 -928 12181 -916
rect 12251 -420 12309 -408
rect 12251 -916 12263 -420
rect 12297 -916 12309 -420
rect 12251 -928 12309 -916
rect 3257 -2945 3457 -2933
rect 3257 -2979 3269 -2945
rect 3445 -2979 3457 -2945
rect 3257 -2991 3457 -2979
rect 3257 -3403 3457 -3391
rect 3257 -3437 3269 -3403
rect 3445 -3437 3457 -3403
rect 3257 -3449 3457 -3437
rect 3257 -3526 3457 -3514
rect 3257 -3560 3269 -3526
rect 3445 -3560 3457 -3526
rect 3257 -3572 3457 -3560
rect 3257 -3984 3457 -3972
rect 3257 -4018 3269 -3984
rect 3445 -4018 3457 -3984
rect 3257 -4030 3457 -4018
rect 3257 -4816 3457 -4804
rect 3257 -4850 3269 -4816
rect 3445 -4850 3457 -4816
rect 3257 -4862 3457 -4850
rect 3257 -5274 3457 -5262
rect 3257 -5308 3269 -5274
rect 3445 -5308 3457 -5274
rect 3257 -5320 3457 -5308
rect 3257 -6106 3457 -6094
rect 3257 -6140 3269 -6106
rect 3445 -6140 3457 -6106
rect 3257 -6152 3457 -6140
rect 3257 -6564 3457 -6552
rect 3257 -6598 3269 -6564
rect 3445 -6598 3457 -6564
rect 3257 -6610 3457 -6598
rect 3257 -7396 3457 -7384
rect 3257 -7430 3269 -7396
rect 3445 -7430 3457 -7396
rect 3257 -7442 3457 -7430
rect 3257 -7854 3457 -7842
rect 3257 -7888 3269 -7854
rect 3445 -7888 3457 -7854
rect 3257 -7900 3457 -7888
rect 3257 -8484 3457 -8472
rect 3257 -8518 3269 -8484
rect 3445 -8518 3457 -8484
rect 3257 -8530 3457 -8518
rect 1926 -9349 2606 -9297
rect 1926 -9383 1978 -9349
rect 2012 -9383 2068 -9349
rect 2102 -9383 2158 -9349
rect 2192 -9383 2248 -9349
rect 2282 -9383 2338 -9349
rect 2372 -9383 2428 -9349
rect 2462 -9383 2518 -9349
rect 2552 -9383 2606 -9349
rect 1926 -9439 2606 -9383
rect 1926 -9473 1978 -9439
rect 2012 -9473 2068 -9439
rect 2102 -9473 2158 -9439
rect 2192 -9473 2248 -9439
rect 2282 -9473 2338 -9439
rect 2372 -9473 2428 -9439
rect 2462 -9473 2518 -9439
rect 2552 -9473 2606 -9439
rect 1926 -9529 2606 -9473
rect 1926 -9563 1978 -9529
rect 2012 -9563 2068 -9529
rect 2102 -9563 2158 -9529
rect 2192 -9563 2248 -9529
rect 2282 -9563 2338 -9529
rect 2372 -9563 2428 -9529
rect 2462 -9563 2518 -9529
rect 2552 -9563 2606 -9529
rect 1926 -9619 2606 -9563
rect 1926 -9653 1978 -9619
rect 2012 -9653 2068 -9619
rect 2102 -9653 2158 -9619
rect 2192 -9653 2248 -9619
rect 2282 -9653 2338 -9619
rect 2372 -9653 2428 -9619
rect 2462 -9653 2518 -9619
rect 2552 -9653 2606 -9619
rect 1926 -9709 2606 -9653
rect 1926 -9743 1978 -9709
rect 2012 -9743 2068 -9709
rect 2102 -9743 2158 -9709
rect 2192 -9743 2248 -9709
rect 2282 -9743 2338 -9709
rect 2372 -9743 2428 -9709
rect 2462 -9743 2518 -9709
rect 2552 -9743 2606 -9709
rect 1926 -9799 2606 -9743
rect 1926 -9833 1978 -9799
rect 2012 -9833 2068 -9799
rect 2102 -9833 2158 -9799
rect 2192 -9833 2248 -9799
rect 2282 -9833 2338 -9799
rect 2372 -9833 2428 -9799
rect 2462 -9833 2518 -9799
rect 2552 -9833 2606 -9799
rect 1926 -9889 2606 -9833
rect 1926 -9923 1978 -9889
rect 2012 -9923 2068 -9889
rect 2102 -9923 2158 -9889
rect 2192 -9923 2248 -9889
rect 2282 -9923 2338 -9889
rect 2372 -9923 2428 -9889
rect 2462 -9923 2518 -9889
rect 2552 -9923 2606 -9889
rect 1926 -9977 2606 -9923
rect 3257 -8742 3457 -8730
rect 3257 -8776 3269 -8742
rect 3445 -8776 3457 -8742
rect 3257 -8788 3457 -8776
rect 3257 -9000 3457 -8988
rect 3257 -9034 3269 -9000
rect 3445 -9034 3457 -9000
rect 3257 -9046 3457 -9034
rect 3257 -9209 3357 -9197
rect 3257 -9243 3269 -9209
rect 3345 -9243 3357 -9209
rect 3257 -9255 3357 -9243
rect 3257 -9667 3357 -9655
rect 3257 -9701 3269 -9667
rect 3345 -9701 3357 -9667
rect 3257 -9713 3357 -9701
rect 3257 -10125 3357 -10113
rect 3257 -10159 3269 -10125
rect 3345 -10159 3357 -10125
rect 3257 -10171 3357 -10159
<< ndiffc >>
rect -10065 1636 -9489 1670
rect -10065 578 -9489 612
rect -8738 2007 -8704 3183
rect -6280 2007 -6246 3183
rect -3822 2007 -3788 3183
rect -8739 132 -8705 1308
rect -6281 132 -6247 1308
rect -3823 132 -3789 1308
rect -1466 -1148 -1432 -872
rect 472 -1148 506 -872
rect 2410 -1148 2444 -872
rect 4348 -1148 4382 -872
rect 6286 -1148 6320 -872
rect -1466 -1558 -1432 -1282
rect 472 -1558 506 -1282
rect 2410 -1558 2444 -1282
rect 4348 -1558 4382 -1282
rect 6286 -1558 6320 -1282
rect 8631 -878 8665 -302
rect 9089 -878 9123 -302
rect 9547 -878 9581 -302
rect 10005 -878 10039 -302
rect 10463 -878 10497 -302
rect 8631 -2085 8665 -1509
rect 9089 -2085 9123 -1509
rect 9547 -2085 9581 -1509
rect 10005 -2085 10039 -1509
rect 10463 -2085 10497 -1509
rect 11819 -1601 11853 -1425
rect 11907 -1601 11941 -1425
rect 12175 -1601 12209 -1425
rect 12263 -1601 12297 -1425
rect -1136 -3849 -360 -3815
rect 345 -3849 1121 -3815
rect -1136 -4107 -360 -4073
rect 345 -4107 1121 -4073
rect -1136 -4365 -360 -4331
rect 345 -4365 1121 -4331
rect -1136 -4623 -360 -4589
rect 345 -4623 1121 -4589
rect -1136 -4881 -360 -4847
rect 345 -4881 1121 -4847
rect -1136 -5139 -360 -5105
rect 345 -5139 1121 -5105
rect -1136 -5397 -360 -5363
rect 345 -5397 1121 -5363
rect -1136 -5655 -360 -5621
rect 345 -5655 1121 -5621
rect -1136 -5913 -360 -5879
rect 345 -5913 1121 -5879
rect -1136 -6171 -360 -6137
rect 345 -6171 1121 -6137
rect -1136 -6429 -360 -6395
rect 345 -6429 1121 -6395
rect -1136 -6687 -360 -6653
rect 345 -6687 1121 -6653
rect -1136 -6945 -360 -6911
rect 345 -6945 1121 -6911
rect -1136 -7203 -360 -7169
rect 345 -7203 1121 -7169
rect -1136 -7461 -360 -7427
rect 345 -7461 1121 -7427
rect -1136 -7719 -360 -7685
rect 345 -7719 1121 -7685
rect -1136 -7977 -360 -7943
rect 345 -7977 1121 -7943
rect -1136 -8235 -360 -8201
rect 345 -8235 1121 -8201
rect -1136 -8493 -360 -8459
rect 345 -8493 1121 -8459
rect -1136 -8751 -360 -8717
rect 345 -8751 1121 -8717
rect -1136 -9009 -360 -8975
rect 345 -9009 1121 -8975
rect -1136 -9267 -360 -9233
rect 345 -9267 1121 -9233
rect -1136 -9525 -360 -9491
rect 345 -9525 1121 -9491
rect -1136 -9783 -360 -9749
rect 345 -9783 1121 -9749
rect -1136 -10041 -360 -10007
rect 345 -10041 1121 -10007
rect 2482 -3044 2658 -3010
rect 2482 -3302 2658 -3268
rect 2482 -3560 2658 -3526
rect 2482 -3818 2658 -3784
rect 2482 -4076 2658 -4042
rect 2482 -4334 2658 -4300
rect 2482 -4592 2658 -4558
rect 2482 -4850 2658 -4816
rect 2482 -5108 2658 -5074
rect 2482 -5366 2658 -5332
rect 2482 -5624 2658 -5590
rect 2482 -5882 2658 -5848
rect 2482 -6140 2658 -6106
rect 2482 -6398 2658 -6364
rect 2482 -6656 2658 -6622
rect 2482 -6914 2658 -6880
rect 2482 -7172 2658 -7138
rect 2482 -7430 2658 -7396
rect 2482 -7688 2658 -7654
rect 2482 -7946 2658 -7912
rect 2482 -8204 2658 -8170
rect 9052 -2669 10128 -2635
rect 9052 -3027 10128 -2993
rect 9052 -3385 10128 -3351
<< pdiffc >>
rect -9948 4719 -9914 5055
rect -6290 4719 -6256 5055
rect -2632 4719 -2598 5055
rect -9948 4231 -9914 4567
rect -6290 4231 -6256 4567
rect -2632 4231 -2598 4567
rect -1476 4155 -1442 7131
rect -1038 4155 -1004 7131
rect -600 4155 -566 7131
rect -162 4155 -128 7131
rect 276 4155 310 7131
rect -1476 178 -1442 3154
rect -1038 178 -1004 3154
rect -600 178 -566 3154
rect -162 178 -128 3154
rect 276 178 310 3154
rect 3353 224 3387 1600
rect 3771 224 3805 1600
rect 4189 224 4223 1600
rect 4607 224 4641 1600
rect 5025 224 5059 1600
rect 7446 1669 7480 2145
rect 8504 1669 8538 2145
rect 9562 1669 9596 2145
rect 10620 1669 10654 2145
rect 11678 1669 11712 2145
rect 7446 507 7480 983
rect 8504 507 8538 983
rect 9562 507 9596 983
rect 10620 507 10654 983
rect 11678 507 11712 983
rect 11779 -916 11813 -420
rect 11907 -916 11941 -420
rect 12135 -916 12169 -420
rect 12263 -916 12297 -420
rect 3269 -2979 3445 -2945
rect 3269 -3437 3445 -3403
rect 3269 -3560 3445 -3526
rect 3269 -4018 3445 -3984
rect 3269 -4850 3445 -4816
rect 3269 -5308 3445 -5274
rect 3269 -6140 3445 -6106
rect 3269 -6598 3445 -6564
rect 3269 -7430 3445 -7396
rect 3269 -7888 3445 -7854
rect 3269 -8518 3445 -8484
rect 1978 -9383 2012 -9349
rect 2068 -9383 2102 -9349
rect 2158 -9383 2192 -9349
rect 2248 -9383 2282 -9349
rect 2338 -9383 2372 -9349
rect 2428 -9383 2462 -9349
rect 2518 -9383 2552 -9349
rect 1978 -9473 2012 -9439
rect 2068 -9473 2102 -9439
rect 2158 -9473 2192 -9439
rect 2248 -9473 2282 -9439
rect 2338 -9473 2372 -9439
rect 2428 -9473 2462 -9439
rect 2518 -9473 2552 -9439
rect 1978 -9563 2012 -9529
rect 2068 -9563 2102 -9529
rect 2158 -9563 2192 -9529
rect 2248 -9563 2282 -9529
rect 2338 -9563 2372 -9529
rect 2428 -9563 2462 -9529
rect 2518 -9563 2552 -9529
rect 1978 -9653 2012 -9619
rect 2068 -9653 2102 -9619
rect 2158 -9653 2192 -9619
rect 2248 -9653 2282 -9619
rect 2338 -9653 2372 -9619
rect 2428 -9653 2462 -9619
rect 2518 -9653 2552 -9619
rect 1978 -9743 2012 -9709
rect 2068 -9743 2102 -9709
rect 2158 -9743 2192 -9709
rect 2248 -9743 2282 -9709
rect 2338 -9743 2372 -9709
rect 2428 -9743 2462 -9709
rect 2518 -9743 2552 -9709
rect 1978 -9833 2012 -9799
rect 2068 -9833 2102 -9799
rect 2158 -9833 2192 -9799
rect 2248 -9833 2282 -9799
rect 2338 -9833 2372 -9799
rect 2428 -9833 2462 -9799
rect 2518 -9833 2552 -9799
rect 1978 -9923 2012 -9889
rect 2068 -9923 2102 -9889
rect 2158 -9923 2192 -9889
rect 2248 -9923 2282 -9889
rect 2338 -9923 2372 -9889
rect 2428 -9923 2462 -9889
rect 2518 -9923 2552 -9889
rect 3269 -8776 3445 -8742
rect 3269 -9034 3445 -9000
rect 3269 -9243 3345 -9209
rect 3269 -9701 3345 -9667
rect 3269 -10159 3345 -10125
<< psubdiff >>
rect -8974 3365 -8914 3399
rect -3613 3365 -3553 3399
rect -8974 3339 -8940 3365
rect -10251 1750 -10155 1784
rect -9399 1750 -9303 1784
rect -10251 1688 -10217 1750
rect -9337 1688 -9303 1750
rect -10251 498 -10217 560
rect -9337 498 -9303 560
rect -10251 464 -10155 498
rect -9399 464 -9303 498
rect -3587 3339 -3553 3365
rect -8974 -29 -8940 -3
rect -3587 -29 -3553 -3
rect -8974 -63 -8914 -29
rect -3613 -63 -3553 -29
rect 8521 -108 8581 -74
rect 10563 -108 10623 -74
rect 8521 -134 8555 -108
rect -1688 -530 -1628 -496
rect 6541 -530 6601 -496
rect -1688 -556 -1654 -530
rect 6567 -556 6601 -530
rect -1688 -1805 -1654 -1779
rect 6567 -1805 6601 -1779
rect -1688 -1839 -1628 -1805
rect 6541 -1839 6601 -1805
rect 10589 -134 10623 -108
rect 8521 -2278 8555 -2252
rect 11697 -1273 11757 -1239
rect 12356 -1273 12416 -1239
rect 11697 -1299 11731 -1273
rect 12382 -1299 12416 -1273
rect 11697 -1765 11731 -1739
rect 12382 -1765 12416 -1739
rect 11697 -1799 11757 -1765
rect 12356 -1799 12416 -1765
rect 10589 -2278 10623 -2252
rect 8521 -2312 8581 -2278
rect 10563 -2312 10623 -2278
rect 11145 -2273 11241 -2239
rect 12381 -2273 12477 -2239
rect 11145 -2335 11179 -2273
rect 12443 -2335 12477 -2273
rect 8866 -2555 8962 -2521
rect 10218 -2555 10314 -2521
rect 8866 -2617 8900 -2555
rect 2224 -2877 2284 -2843
rect 2866 -2877 2926 -2843
rect 2224 -2903 2258 -2877
rect -1424 -3705 -1364 -3671
rect 1345 -3705 1405 -3671
rect -1424 -3731 -1390 -3705
rect 1371 -3731 1405 -3705
rect -1424 -10213 -1390 -10187
rect 2892 -2903 2926 -2877
rect 2224 -8337 2258 -8311
rect 10280 -2617 10314 -2555
rect 11145 -2535 11179 -2473
rect 12443 -2535 12477 -2473
rect 11145 -2569 11241 -2535
rect 12381 -2569 12477 -2535
rect 8866 -3465 8900 -3403
rect 10280 -3465 10314 -3403
rect 8866 -3499 8962 -3465
rect 10218 -3499 10314 -3465
rect 2892 -8337 2926 -8311
rect 2224 -8371 2284 -8337
rect 2866 -8371 2926 -8337
rect 1371 -10213 1405 -10187
rect -1424 -10247 -1364 -10213
rect 1345 -10247 1405 -10213
rect 1622 -9026 2910 -8993
rect 1622 -9060 1680 -9026
rect 1714 -9060 1770 -9026
rect 1804 -9060 1860 -9026
rect 1894 -9060 1950 -9026
rect 1984 -9060 2040 -9026
rect 2074 -9060 2130 -9026
rect 2164 -9060 2220 -9026
rect 2254 -9060 2310 -9026
rect 2344 -9060 2400 -9026
rect 2434 -9060 2490 -9026
rect 2524 -9060 2580 -9026
rect 2614 -9060 2670 -9026
rect 2704 -9060 2760 -9026
rect 2794 -9060 2910 -9026
rect 1622 -9094 2910 -9060
rect 1622 -9127 1723 -9094
rect 1622 -9161 1657 -9127
rect 1691 -9161 1723 -9127
rect 2809 -9127 2910 -9094
rect 1622 -9217 1723 -9161
rect 1622 -9251 1657 -9217
rect 1691 -9251 1723 -9217
rect 1622 -9307 1723 -9251
rect 1622 -9341 1657 -9307
rect 1691 -9341 1723 -9307
rect 1622 -9397 1723 -9341
rect 1622 -9431 1657 -9397
rect 1691 -9431 1723 -9397
rect 1622 -9487 1723 -9431
rect 1622 -9521 1657 -9487
rect 1691 -9521 1723 -9487
rect 1622 -9577 1723 -9521
rect 1622 -9611 1657 -9577
rect 1691 -9611 1723 -9577
rect 1622 -9667 1723 -9611
rect 1622 -9701 1657 -9667
rect 1691 -9701 1723 -9667
rect 1622 -9757 1723 -9701
rect 1622 -9791 1657 -9757
rect 1691 -9791 1723 -9757
rect 1622 -9847 1723 -9791
rect 1622 -9881 1657 -9847
rect 1691 -9881 1723 -9847
rect 1622 -9937 1723 -9881
rect 1622 -9971 1657 -9937
rect 1691 -9971 1723 -9937
rect 1622 -10027 1723 -9971
rect 1622 -10061 1657 -10027
rect 1691 -10061 1723 -10027
rect 1622 -10117 1723 -10061
rect 1622 -10151 1657 -10117
rect 1691 -10151 1723 -10117
rect 2809 -9161 2844 -9127
rect 2878 -9161 2910 -9127
rect 2809 -9217 2910 -9161
rect 2809 -9251 2844 -9217
rect 2878 -9251 2910 -9217
rect 2809 -9307 2910 -9251
rect 2809 -9341 2844 -9307
rect 2878 -9341 2910 -9307
rect 2809 -9397 2910 -9341
rect 2809 -9431 2844 -9397
rect 2878 -9431 2910 -9397
rect 2809 -9487 2910 -9431
rect 2809 -9521 2844 -9487
rect 2878 -9521 2910 -9487
rect 2809 -9577 2910 -9521
rect 2809 -9611 2844 -9577
rect 2878 -9611 2910 -9577
rect 2809 -9667 2910 -9611
rect 2809 -9701 2844 -9667
rect 2878 -9701 2910 -9667
rect 2809 -9757 2910 -9701
rect 2809 -9791 2844 -9757
rect 2878 -9791 2910 -9757
rect 2809 -9847 2910 -9791
rect 2809 -9881 2844 -9847
rect 2878 -9881 2910 -9847
rect 2809 -9937 2910 -9881
rect 2809 -9971 2844 -9937
rect 2878 -9971 2910 -9937
rect 2809 -10027 2910 -9971
rect 2809 -10061 2844 -10027
rect 2878 -10061 2910 -10027
rect 2809 -10117 2910 -10061
rect 1622 -10180 1723 -10151
rect 2809 -10151 2844 -10117
rect 2878 -10151 2910 -10117
rect 2809 -10180 2910 -10151
rect 1622 -10213 2910 -10180
rect 1622 -10247 1680 -10213
rect 1714 -10247 1770 -10213
rect 1804 -10247 1860 -10213
rect 1894 -10247 1950 -10213
rect 1984 -10247 2040 -10213
rect 2074 -10247 2130 -10213
rect 2164 -10247 2220 -10213
rect 2254 -10247 2310 -10213
rect 2344 -10247 2400 -10213
rect 2434 -10247 2490 -10213
rect 2524 -10247 2580 -10213
rect 2614 -10247 2670 -10213
rect 2704 -10247 2760 -10213
rect 2794 -10247 2910 -10213
rect 1622 -10281 2910 -10247
<< nsubdiff >>
rect -1740 7523 -1680 7557
rect 600 7523 660 7557
rect -1740 7497 -1706 7523
rect -10205 5326 -10145 5360
rect -2457 5326 -2397 5360
rect -10205 5300 -10171 5326
rect -2431 5300 -2397 5326
rect -10205 4018 -10171 4044
rect -2431 4018 -2397 4044
rect -10205 3984 -10145 4018
rect -2457 3984 -2397 4018
rect 626 7497 660 7523
rect -1740 -64 -1706 -38
rect 7181 2439 7241 2473
rect 11927 2439 11987 2473
rect 7181 2413 7215 2439
rect 3239 1761 3335 1795
rect 5077 1761 5173 1795
rect 3239 1699 3273 1761
rect 5139 1699 5173 1761
rect 3239 63 3273 125
rect 11953 2413 11987 2439
rect 7181 174 7215 200
rect 11953 174 11987 200
rect 7181 140 7241 174
rect 11927 140 11987 174
rect 5139 63 5173 125
rect 3239 29 3335 63
rect 5077 29 5173 63
rect 626 -64 660 -38
rect -1740 -98 -1680 -64
rect 600 -98 660 -64
rect 11665 -259 11761 -225
rect 11959 -259 12117 -225
rect 12315 -259 12411 -225
rect 11665 -321 11699 -259
rect 12021 -321 12055 -259
rect 11665 -1077 11699 -1015
rect 12377 -321 12411 -259
rect 12021 -1077 12055 -1015
rect 12377 -1077 12411 -1015
rect 11665 -1111 11761 -1077
rect 11959 -1111 12117 -1077
rect 12315 -1111 12411 -1077
rect 3098 -2869 3158 -2835
rect 3582 -2869 3642 -2835
rect 3098 -2895 3132 -2869
rect 3608 -2895 3642 -2869
rect 3098 -4085 3132 -4059
rect 3608 -4085 3642 -4059
rect 3098 -4119 3158 -4085
rect 3582 -4119 3642 -4085
rect 3074 -4736 3170 -4702
rect 3544 -4736 3640 -4702
rect 3074 -4798 3108 -4736
rect 3606 -4798 3640 -4736
rect 3074 -5388 3108 -5326
rect 3606 -5388 3640 -5326
rect 3074 -5422 3170 -5388
rect 3544 -5422 3640 -5388
rect 3074 -6026 3170 -5992
rect 3544 -6026 3640 -5992
rect 3074 -6088 3108 -6026
rect 3606 -6088 3640 -6026
rect 3074 -6678 3108 -6616
rect 3606 -6678 3640 -6616
rect 3074 -6712 3170 -6678
rect 3544 -6712 3640 -6678
rect 3074 -7316 3170 -7282
rect 3544 -7316 3640 -7282
rect 3074 -7378 3108 -7316
rect 3606 -7378 3640 -7316
rect 3074 -7968 3108 -7906
rect 3606 -7968 3640 -7906
rect 3074 -8002 3170 -7968
rect 3544 -8002 3640 -7968
rect 3083 -8417 3166 -8368
rect 3545 -8417 3633 -8368
rect 3083 -8479 3131 -8417
rect 3581 -8486 3633 -8417
rect 1785 -9175 2747 -9156
rect 1785 -9209 1880 -9175
rect 1914 -9209 1970 -9175
rect 2004 -9209 2060 -9175
rect 2094 -9209 2150 -9175
rect 2184 -9209 2240 -9175
rect 2274 -9209 2330 -9175
rect 2364 -9209 2420 -9175
rect 2454 -9209 2510 -9175
rect 2544 -9209 2600 -9175
rect 2634 -9209 2747 -9175
rect 1785 -9228 2747 -9209
rect 1785 -9233 1857 -9228
rect 1785 -9267 1804 -9233
rect 1838 -9267 1857 -9233
rect 1785 -9323 1857 -9267
rect 2675 -9267 2747 -9228
rect 1785 -9357 1804 -9323
rect 1838 -9357 1857 -9323
rect 1785 -9413 1857 -9357
rect 1785 -9447 1804 -9413
rect 1838 -9447 1857 -9413
rect 1785 -9503 1857 -9447
rect 1785 -9537 1804 -9503
rect 1838 -9537 1857 -9503
rect 1785 -9593 1857 -9537
rect 1785 -9627 1804 -9593
rect 1838 -9627 1857 -9593
rect 1785 -9683 1857 -9627
rect 1785 -9717 1804 -9683
rect 1838 -9717 1857 -9683
rect 1785 -9773 1857 -9717
rect 1785 -9807 1804 -9773
rect 1838 -9807 1857 -9773
rect 1785 -9863 1857 -9807
rect 1785 -9897 1804 -9863
rect 1838 -9897 1857 -9863
rect 1785 -9953 1857 -9897
rect 1785 -9987 1804 -9953
rect 1838 -9987 1857 -9953
rect 2675 -9301 2694 -9267
rect 2728 -9301 2747 -9267
rect 2675 -9357 2747 -9301
rect 2675 -9391 2694 -9357
rect 2728 -9391 2747 -9357
rect 2675 -9447 2747 -9391
rect 2675 -9481 2694 -9447
rect 2728 -9481 2747 -9447
rect 2675 -9537 2747 -9481
rect 2675 -9571 2694 -9537
rect 2728 -9571 2747 -9537
rect 2675 -9627 2747 -9571
rect 2675 -9661 2694 -9627
rect 2728 -9661 2747 -9627
rect 2675 -9717 2747 -9661
rect 2675 -9751 2694 -9717
rect 2728 -9751 2747 -9717
rect 2675 -9807 2747 -9751
rect 2675 -9841 2694 -9807
rect 2728 -9841 2747 -9807
rect 2675 -9897 2747 -9841
rect 2675 -9931 2694 -9897
rect 2728 -9931 2747 -9897
rect 1785 -10046 1857 -9987
rect 2675 -9987 2747 -9931
rect 2675 -10021 2694 -9987
rect 2728 -10021 2747 -9987
rect 2675 -10046 2747 -10021
rect 1785 -10065 2747 -10046
rect 1785 -10099 1861 -10065
rect 1895 -10099 1951 -10065
rect 1985 -10099 2041 -10065
rect 2075 -10099 2131 -10065
rect 2165 -10099 2221 -10065
rect 2255 -10099 2311 -10065
rect 2345 -10099 2401 -10065
rect 2435 -10099 2491 -10065
rect 2525 -10099 2581 -10065
rect 2615 -10099 2747 -10065
rect 1785 -10118 2747 -10099
rect 3083 -9013 3131 -8756
rect 3083 -10257 3131 -10121
rect 3581 -10257 3633 -10161
rect 3083 -10309 3250 -10257
rect 3486 -10309 3633 -10257
<< psubdiffcont >>
rect -8914 3365 -3613 3399
rect -10155 1750 -9399 1784
rect -10251 560 -10217 1688
rect -9337 560 -9303 1688
rect -10155 464 -9399 498
rect -8974 -3 -8940 3339
rect -3587 -3 -3553 3339
rect -8914 -63 -3613 -29
rect 8581 -108 10563 -74
rect -1628 -530 6541 -496
rect -1688 -1779 -1654 -556
rect 6567 -1779 6601 -556
rect -1628 -1839 6541 -1805
rect 8521 -2252 8555 -134
rect 10589 -2252 10623 -134
rect 11757 -1273 12356 -1239
rect 11697 -1739 11731 -1299
rect 12382 -1739 12416 -1299
rect 11757 -1799 12356 -1765
rect 8581 -2312 10563 -2278
rect 11241 -2273 12381 -2239
rect 11145 -2473 11179 -2335
rect 8962 -2555 10218 -2521
rect 2284 -2877 2866 -2843
rect -1364 -3705 1345 -3671
rect -1424 -10187 -1390 -3731
rect 1371 -10187 1405 -3731
rect 2224 -8311 2258 -2903
rect 2892 -8311 2926 -2903
rect 8866 -3403 8900 -2617
rect 12443 -2473 12477 -2335
rect 11241 -2569 12381 -2535
rect 10280 -3403 10314 -2617
rect 8962 -3499 10218 -3465
rect 2284 -8371 2866 -8337
rect -1364 -10247 1345 -10213
rect 1680 -9060 1714 -9026
rect 1770 -9060 1804 -9026
rect 1860 -9060 1894 -9026
rect 1950 -9060 1984 -9026
rect 2040 -9060 2074 -9026
rect 2130 -9060 2164 -9026
rect 2220 -9060 2254 -9026
rect 2310 -9060 2344 -9026
rect 2400 -9060 2434 -9026
rect 2490 -9060 2524 -9026
rect 2580 -9060 2614 -9026
rect 2670 -9060 2704 -9026
rect 2760 -9060 2794 -9026
rect 1657 -9161 1691 -9127
rect 1657 -9251 1691 -9217
rect 1657 -9341 1691 -9307
rect 1657 -9431 1691 -9397
rect 1657 -9521 1691 -9487
rect 1657 -9611 1691 -9577
rect 1657 -9701 1691 -9667
rect 1657 -9791 1691 -9757
rect 1657 -9881 1691 -9847
rect 1657 -9971 1691 -9937
rect 1657 -10061 1691 -10027
rect 1657 -10151 1691 -10117
rect 2844 -9161 2878 -9127
rect 2844 -9251 2878 -9217
rect 2844 -9341 2878 -9307
rect 2844 -9431 2878 -9397
rect 2844 -9521 2878 -9487
rect 2844 -9611 2878 -9577
rect 2844 -9701 2878 -9667
rect 2844 -9791 2878 -9757
rect 2844 -9881 2878 -9847
rect 2844 -9971 2878 -9937
rect 2844 -10061 2878 -10027
rect 2844 -10151 2878 -10117
rect 1680 -10247 1714 -10213
rect 1770 -10247 1804 -10213
rect 1860 -10247 1894 -10213
rect 1950 -10247 1984 -10213
rect 2040 -10247 2074 -10213
rect 2130 -10247 2164 -10213
rect 2220 -10247 2254 -10213
rect 2310 -10247 2344 -10213
rect 2400 -10247 2434 -10213
rect 2490 -10247 2524 -10213
rect 2580 -10247 2614 -10213
rect 2670 -10247 2704 -10213
rect 2760 -10247 2794 -10213
<< nsubdiffcont >>
rect -1680 7523 600 7557
rect -10145 5326 -2457 5360
rect -10205 4044 -10171 5300
rect -2431 4044 -2397 5300
rect -10145 3984 -2457 4018
rect -1740 -38 -1706 7497
rect 626 -38 660 7497
rect 7241 2439 11927 2473
rect 3335 1761 5077 1795
rect 3239 125 3273 1699
rect 5139 125 5173 1699
rect 7181 200 7215 2413
rect 11953 200 11987 2413
rect 7241 140 11927 174
rect 3335 29 5077 63
rect -1680 -98 600 -64
rect 11761 -259 11959 -225
rect 12117 -259 12315 -225
rect 11665 -1015 11699 -321
rect 12021 -1015 12055 -321
rect 12377 -1015 12411 -321
rect 11761 -1111 11959 -1077
rect 12117 -1111 12315 -1077
rect 3158 -2869 3582 -2835
rect 3098 -4059 3132 -2895
rect 3608 -4059 3642 -2895
rect 3158 -4119 3582 -4085
rect 3170 -4736 3544 -4702
rect 3074 -5326 3108 -4798
rect 3606 -5326 3640 -4798
rect 3170 -5422 3544 -5388
rect 3170 -6026 3544 -5992
rect 3074 -6616 3108 -6088
rect 3606 -6616 3640 -6088
rect 3170 -6712 3544 -6678
rect 3170 -7316 3544 -7282
rect 3074 -7906 3108 -7378
rect 3606 -7906 3640 -7378
rect 3170 -8002 3544 -7968
rect 3166 -8417 3545 -8368
rect 3083 -8756 3131 -8479
rect 1880 -9209 1914 -9175
rect 1970 -9209 2004 -9175
rect 2060 -9209 2094 -9175
rect 2150 -9209 2184 -9175
rect 2240 -9209 2274 -9175
rect 2330 -9209 2364 -9175
rect 2420 -9209 2454 -9175
rect 2510 -9209 2544 -9175
rect 2600 -9209 2634 -9175
rect 1804 -9267 1838 -9233
rect 1804 -9357 1838 -9323
rect 1804 -9447 1838 -9413
rect 1804 -9537 1838 -9503
rect 1804 -9627 1838 -9593
rect 1804 -9717 1838 -9683
rect 1804 -9807 1838 -9773
rect 1804 -9897 1838 -9863
rect 1804 -9987 1838 -9953
rect 2694 -9301 2728 -9267
rect 2694 -9391 2728 -9357
rect 2694 -9481 2728 -9447
rect 2694 -9571 2728 -9537
rect 2694 -9661 2728 -9627
rect 2694 -9751 2728 -9717
rect 2694 -9841 2728 -9807
rect 2694 -9931 2728 -9897
rect 2694 -10021 2728 -9987
rect 1861 -10099 1895 -10065
rect 1951 -10099 1985 -10065
rect 2041 -10099 2075 -10065
rect 2131 -10099 2165 -10065
rect 2221 -10099 2255 -10065
rect 2311 -10099 2345 -10065
rect 2401 -10099 2435 -10065
rect 2491 -10099 2525 -10065
rect 2581 -10099 2615 -10065
rect 3083 -10121 3131 -9013
rect 3581 -10161 3633 -8486
rect 3250 -10309 3486 -10257
<< poly >>
rect -9902 5148 -6302 5164
rect -9902 5114 -9886 5148
rect -6318 5114 -6302 5148
rect -9902 5067 -6302 5114
rect -6244 5148 -2644 5164
rect -6244 5114 -6228 5148
rect -2660 5114 -2644 5148
rect -6244 5067 -2644 5114
rect -9902 4660 -6302 4707
rect -9902 4626 -9886 4660
rect -6318 4626 -6302 4660
rect -9902 4579 -6302 4626
rect -6244 4660 -2644 4707
rect -6244 4626 -6228 4660
rect -2660 4626 -2644 4660
rect -6244 4579 -2644 4626
rect -9902 4172 -6302 4219
rect -9902 4138 -9886 4172
rect -6318 4138 -6302 4172
rect -9902 4122 -6302 4138
rect -6244 4172 -2644 4219
rect -6244 4138 -6228 4172
rect -2660 4138 -2644 4172
rect -6244 4122 -2644 4138
rect -10165 1608 -10077 1624
rect -10165 640 -10149 1608
rect -10115 640 -10077 1608
rect -10165 624 -10077 640
rect -9477 1608 -9389 1624
rect -9477 640 -9439 1608
rect -9405 640 -9389 1608
rect -9477 624 -9389 640
rect -8692 3267 -6292 3283
rect -8692 3233 -8676 3267
rect -6308 3233 -6292 3267
rect -8692 3195 -6292 3233
rect -6234 3267 -3834 3283
rect -6234 3233 -6218 3267
rect -3850 3233 -3834 3267
rect -6234 3195 -3834 3233
rect -8692 1957 -6292 1995
rect -8692 1923 -8676 1957
rect -6308 1923 -6292 1957
rect -8692 1907 -6292 1923
rect -6234 1957 -3834 1995
rect -6234 1923 -6218 1957
rect -3850 1923 -3834 1957
rect -6234 1907 -3834 1923
rect -8693 1392 -6293 1408
rect -8693 1358 -8677 1392
rect -6309 1358 -6293 1392
rect -8693 1320 -6293 1358
rect -6235 1392 -3835 1408
rect -6235 1358 -6219 1392
rect -3851 1358 -3835 1392
rect -6235 1320 -3835 1358
rect -8693 82 -6293 120
rect -8693 48 -8677 82
rect -6309 48 -6293 82
rect -8693 32 -6293 48
rect -6235 82 -3835 120
rect -6235 48 -6219 82
rect -3851 48 -3835 82
rect -6235 32 -3835 48
rect -1430 7224 -1050 7240
rect -1430 7190 -1414 7224
rect -1066 7190 -1050 7224
rect -1430 7143 -1050 7190
rect -992 7224 -612 7240
rect -992 7190 -976 7224
rect -628 7190 -612 7224
rect -992 7143 -612 7190
rect -554 7224 -174 7240
rect -554 7190 -538 7224
rect -190 7190 -174 7224
rect -554 7143 -174 7190
rect -116 7224 264 7240
rect -116 7190 -100 7224
rect 248 7190 264 7224
rect -116 7143 264 7190
rect -1430 4096 -1050 4143
rect -1430 4062 -1414 4096
rect -1066 4062 -1050 4096
rect -1430 4046 -1050 4062
rect -992 4096 -612 4143
rect -992 4062 -976 4096
rect -628 4062 -612 4096
rect -992 4046 -612 4062
rect -554 4096 -174 4143
rect -554 4062 -538 4096
rect -190 4062 -174 4096
rect -554 4046 -174 4062
rect -116 4096 264 4143
rect -116 4062 -100 4096
rect 248 4062 264 4096
rect -116 4046 264 4062
rect -1430 3247 -1050 3263
rect -1430 3213 -1414 3247
rect -1066 3213 -1050 3247
rect -1430 3166 -1050 3213
rect -992 3247 -612 3263
rect -992 3213 -976 3247
rect -628 3213 -612 3247
rect -992 3166 -612 3213
rect -554 3247 -174 3263
rect -554 3213 -538 3247
rect -190 3213 -174 3247
rect -554 3166 -174 3213
rect -116 3247 264 3263
rect -116 3213 -100 3247
rect 248 3213 264 3247
rect -116 3166 264 3213
rect -1430 119 -1050 166
rect -1430 85 -1414 119
rect -1066 85 -1050 119
rect -1430 69 -1050 85
rect -992 119 -612 166
rect -992 85 -976 119
rect -628 85 -612 119
rect -992 69 -612 85
rect -554 119 -174 166
rect -554 85 -538 119
rect -190 85 -174 119
rect -554 69 -174 85
rect -116 119 264 166
rect -116 85 -100 119
rect 248 85 264 119
rect -116 69 264 85
rect 3399 1693 3759 1709
rect 3399 1659 3415 1693
rect 3743 1659 3759 1693
rect 3399 1612 3759 1659
rect 3817 1693 4177 1709
rect 3817 1659 3833 1693
rect 4161 1659 4177 1693
rect 3817 1612 4177 1659
rect 4235 1693 4595 1709
rect 4235 1659 4251 1693
rect 4579 1659 4595 1693
rect 4235 1612 4595 1659
rect 4653 1693 5013 1709
rect 4653 1659 4669 1693
rect 4997 1659 5013 1693
rect 4653 1612 5013 1659
rect 3399 165 3759 212
rect 3399 131 3415 165
rect 3743 131 3759 165
rect 3399 115 3759 131
rect 3817 165 4177 212
rect 3817 131 3833 165
rect 4161 131 4177 165
rect 3817 115 4177 131
rect 4235 165 4595 212
rect 4235 131 4251 165
rect 4579 131 4595 165
rect 4235 115 4595 131
rect 4653 165 5013 212
rect 4653 131 4669 165
rect 4997 131 5013 165
rect 4653 115 5013 131
rect 7492 2238 8492 2254
rect 7492 2204 7508 2238
rect 8476 2204 8492 2238
rect 7492 2157 8492 2204
rect 8550 2238 9550 2254
rect 8550 2204 8566 2238
rect 9534 2204 9550 2238
rect 8550 2157 9550 2204
rect 9608 2238 10608 2254
rect 9608 2204 9624 2238
rect 10592 2204 10608 2238
rect 9608 2157 10608 2204
rect 10666 2238 11666 2254
rect 10666 2204 10682 2238
rect 11650 2204 11666 2238
rect 10666 2157 11666 2204
rect 7492 1610 8492 1657
rect 7492 1576 7508 1610
rect 8476 1576 8492 1610
rect 7492 1560 8492 1576
rect 8550 1610 9550 1657
rect 8550 1576 8566 1610
rect 9534 1576 9550 1610
rect 8550 1560 9550 1576
rect 9608 1610 10608 1657
rect 9608 1576 9624 1610
rect 10592 1576 10608 1610
rect 9608 1560 10608 1576
rect 10666 1610 11666 1657
rect 10666 1576 10682 1610
rect 11650 1576 11666 1610
rect 10666 1560 11666 1576
rect 7492 1076 8492 1092
rect 7492 1042 7508 1076
rect 8476 1042 8492 1076
rect 7492 995 8492 1042
rect 8550 1076 9550 1092
rect 8550 1042 8566 1076
rect 9534 1042 9550 1076
rect 8550 995 9550 1042
rect 9608 1076 10608 1092
rect 9608 1042 9624 1076
rect 10592 1042 10608 1076
rect 9608 995 10608 1042
rect 10666 1076 11666 1092
rect 10666 1042 10682 1076
rect 11650 1042 11666 1076
rect 10666 995 11666 1042
rect 7492 448 8492 495
rect 7492 414 7508 448
rect 8476 414 8492 448
rect 7492 398 8492 414
rect 8550 448 9550 495
rect 8550 414 8566 448
rect 9534 414 9550 448
rect 8550 398 9550 414
rect 9608 448 10608 495
rect 9608 414 9624 448
rect 10592 414 10608 448
rect 9608 398 10608 414
rect 10666 448 11666 495
rect 10666 414 10682 448
rect 11650 414 11666 448
rect 10666 398 11666 414
rect -1420 -788 460 -772
rect -1420 -822 -1404 -788
rect 444 -822 460 -788
rect -1420 -860 460 -822
rect 518 -788 2398 -772
rect 518 -822 534 -788
rect 2382 -822 2398 -788
rect 518 -860 2398 -822
rect 2456 -788 4336 -772
rect 2456 -822 2472 -788
rect 4320 -822 4336 -788
rect 2456 -860 4336 -822
rect 4394 -788 6274 -772
rect 4394 -822 4410 -788
rect 6258 -822 6274 -788
rect 4394 -860 6274 -822
rect -1420 -1198 460 -1160
rect -1420 -1232 -1404 -1198
rect 444 -1232 460 -1198
rect -1420 -1270 460 -1232
rect 518 -1198 2398 -1160
rect 518 -1232 534 -1198
rect 2382 -1232 2398 -1198
rect 518 -1270 2398 -1232
rect 2456 -1198 4336 -1160
rect 2456 -1232 2472 -1198
rect 4320 -1232 4336 -1198
rect 2456 -1270 4336 -1232
rect 4394 -1198 6274 -1160
rect 4394 -1232 4410 -1198
rect 6258 -1232 6274 -1198
rect 4394 -1270 6274 -1232
rect -1420 -1608 460 -1570
rect -1420 -1642 -1404 -1608
rect 444 -1642 460 -1608
rect -1420 -1658 460 -1642
rect 518 -1608 2398 -1570
rect 518 -1642 534 -1608
rect 2382 -1642 2398 -1608
rect 518 -1658 2398 -1642
rect 2456 -1608 4336 -1570
rect 2456 -1642 2472 -1608
rect 4320 -1642 4336 -1608
rect 2456 -1658 4336 -1642
rect 4394 -1608 6274 -1570
rect 4394 -1642 4410 -1608
rect 6258 -1642 6274 -1608
rect 4394 -1658 6274 -1642
rect 8677 -218 9077 -202
rect 8677 -252 8693 -218
rect 9061 -252 9077 -218
rect 8677 -290 9077 -252
rect 9135 -218 9535 -202
rect 9135 -252 9151 -218
rect 9519 -252 9535 -218
rect 9135 -290 9535 -252
rect 9593 -218 9993 -202
rect 9593 -252 9609 -218
rect 9977 -252 9993 -218
rect 9593 -290 9993 -252
rect 10051 -218 10451 -202
rect 10051 -252 10067 -218
rect 10435 -252 10451 -218
rect 10051 -290 10451 -252
rect 8677 -928 9077 -890
rect 8677 -962 8693 -928
rect 9061 -962 9077 -928
rect 8677 -978 9077 -962
rect 9135 -928 9535 -890
rect 9135 -962 9151 -928
rect 9519 -962 9535 -928
rect 9135 -978 9535 -962
rect 9593 -928 9993 -890
rect 9593 -962 9609 -928
rect 9977 -962 9993 -928
rect 9593 -978 9993 -962
rect 10051 -928 10451 -890
rect 10051 -962 10067 -928
rect 10435 -962 10451 -928
rect 10051 -978 10451 -962
rect 8677 -1425 9077 -1409
rect 8677 -1459 8693 -1425
rect 9061 -1459 9077 -1425
rect 8677 -1497 9077 -1459
rect 9135 -1425 9535 -1409
rect 9135 -1459 9151 -1425
rect 9519 -1459 9535 -1425
rect 9135 -1497 9535 -1459
rect 9593 -1425 9993 -1409
rect 9593 -1459 9609 -1425
rect 9977 -1459 9993 -1425
rect 9593 -1497 9993 -1459
rect 10051 -1425 10451 -1409
rect 10051 -1459 10067 -1425
rect 10435 -1459 10451 -1425
rect 10051 -1497 10451 -1459
rect 8677 -2135 9077 -2097
rect 8677 -2169 8693 -2135
rect 9061 -2169 9077 -2135
rect 8677 -2185 9077 -2169
rect 9135 -2135 9535 -2097
rect 9135 -2169 9151 -2135
rect 9519 -2169 9535 -2135
rect 9135 -2185 9535 -2169
rect 9593 -2135 9993 -2097
rect 9593 -2169 9609 -2135
rect 9977 -2169 9993 -2135
rect 9593 -2185 9993 -2169
rect 10051 -2135 10451 -2097
rect 10051 -2169 10067 -2135
rect 10435 -2169 10451 -2135
rect 10051 -2185 10451 -2169
rect 11825 -327 11895 -311
rect 11825 -361 11841 -327
rect 11879 -361 11895 -327
rect 11825 -408 11895 -361
rect 11825 -975 11895 -928
rect 11825 -1009 11841 -975
rect 11879 -1009 11895 -975
rect 11825 -1025 11895 -1009
rect 12181 -327 12251 -311
rect 12181 -361 12197 -327
rect 12235 -361 12251 -327
rect 12181 -408 12251 -361
rect 12181 -975 12251 -928
rect 12181 -1009 12197 -975
rect 12235 -1009 12251 -975
rect 12181 -1025 12251 -1009
rect 11847 -1341 11913 -1325
rect 11847 -1375 11863 -1341
rect 11897 -1375 11913 -1341
rect 11847 -1391 11913 -1375
rect 12203 -1341 12269 -1325
rect 12203 -1375 12219 -1341
rect 12253 -1375 12269 -1341
rect 12203 -1391 12269 -1375
rect 11865 -1413 11895 -1391
rect 12221 -1413 12251 -1391
rect 11865 -1635 11895 -1613
rect 12221 -1635 12251 -1613
rect 11847 -1651 11913 -1635
rect 11847 -1685 11863 -1651
rect 11897 -1685 11913 -1651
rect 11847 -1701 11913 -1685
rect 12203 -1651 12269 -1635
rect 12203 -1685 12219 -1651
rect 12253 -1685 12269 -1651
rect 12203 -1701 12269 -1685
rect -1236 -3877 -1148 -3861
rect -1236 -4045 -1220 -3877
rect -1186 -4045 -1148 -3877
rect -1236 -4061 -1148 -4045
rect -348 -3877 -260 -3861
rect -348 -4045 -310 -3877
rect -276 -4045 -260 -3877
rect -348 -4061 -260 -4045
rect 245 -3877 333 -3861
rect 245 -4045 261 -3877
rect 295 -4045 333 -3877
rect 245 -4061 333 -4045
rect 1133 -3877 1221 -3861
rect 1133 -4045 1171 -3877
rect 1205 -4045 1221 -3877
rect 1133 -4061 1221 -4045
rect -1236 -4135 -1148 -4119
rect -1236 -4303 -1220 -4135
rect -1186 -4303 -1148 -4135
rect -1236 -4319 -1148 -4303
rect -348 -4135 -260 -4119
rect -348 -4303 -310 -4135
rect -276 -4303 -260 -4135
rect -348 -4319 -260 -4303
rect 245 -4135 333 -4119
rect 245 -4303 261 -4135
rect 295 -4303 333 -4135
rect 245 -4319 333 -4303
rect 1133 -4135 1221 -4119
rect 1133 -4303 1171 -4135
rect 1205 -4303 1221 -4135
rect 1133 -4319 1221 -4303
rect -1236 -4393 -1148 -4377
rect -1236 -4561 -1220 -4393
rect -1186 -4561 -1148 -4393
rect -1236 -4577 -1148 -4561
rect -348 -4393 -260 -4377
rect -348 -4561 -310 -4393
rect -276 -4561 -260 -4393
rect -348 -4577 -260 -4561
rect 245 -4393 333 -4377
rect 245 -4561 261 -4393
rect 295 -4561 333 -4393
rect 245 -4577 333 -4561
rect 1133 -4393 1221 -4377
rect 1133 -4561 1171 -4393
rect 1205 -4561 1221 -4393
rect 1133 -4577 1221 -4561
rect -1236 -4651 -1148 -4635
rect -1236 -4819 -1220 -4651
rect -1186 -4819 -1148 -4651
rect -1236 -4835 -1148 -4819
rect -348 -4651 -260 -4635
rect -348 -4819 -310 -4651
rect -276 -4819 -260 -4651
rect -348 -4835 -260 -4819
rect 245 -4651 333 -4635
rect 245 -4819 261 -4651
rect 295 -4819 333 -4651
rect 245 -4835 333 -4819
rect 1133 -4651 1221 -4635
rect 1133 -4819 1171 -4651
rect 1205 -4819 1221 -4651
rect 1133 -4835 1221 -4819
rect -1236 -4909 -1148 -4893
rect -1236 -5077 -1220 -4909
rect -1186 -5077 -1148 -4909
rect -1236 -5093 -1148 -5077
rect -348 -4909 -260 -4893
rect -348 -5077 -310 -4909
rect -276 -5077 -260 -4909
rect -348 -5093 -260 -5077
rect 245 -4909 333 -4893
rect 245 -5077 261 -4909
rect 295 -5077 333 -4909
rect 245 -5093 333 -5077
rect 1133 -4909 1221 -4893
rect 1133 -5077 1171 -4909
rect 1205 -5077 1221 -4909
rect 1133 -5093 1221 -5077
rect -1236 -5167 -1148 -5151
rect -1236 -5335 -1220 -5167
rect -1186 -5335 -1148 -5167
rect -1236 -5351 -1148 -5335
rect -348 -5167 -260 -5151
rect -348 -5335 -310 -5167
rect -276 -5335 -260 -5167
rect -348 -5351 -260 -5335
rect 245 -5167 333 -5151
rect 245 -5335 261 -5167
rect 295 -5335 333 -5167
rect 245 -5351 333 -5335
rect 1133 -5167 1221 -5151
rect 1133 -5335 1171 -5167
rect 1205 -5335 1221 -5167
rect 1133 -5351 1221 -5335
rect -1236 -5425 -1148 -5409
rect -1236 -5593 -1220 -5425
rect -1186 -5593 -1148 -5425
rect -1236 -5609 -1148 -5593
rect -348 -5425 -260 -5409
rect -348 -5593 -310 -5425
rect -276 -5593 -260 -5425
rect -348 -5609 -260 -5593
rect 245 -5425 333 -5409
rect 245 -5593 261 -5425
rect 295 -5593 333 -5425
rect 245 -5609 333 -5593
rect 1133 -5425 1221 -5409
rect 1133 -5593 1171 -5425
rect 1205 -5593 1221 -5425
rect 1133 -5609 1221 -5593
rect -1236 -5683 -1148 -5667
rect -1236 -5851 -1220 -5683
rect -1186 -5851 -1148 -5683
rect -1236 -5867 -1148 -5851
rect -348 -5683 -260 -5667
rect -348 -5851 -310 -5683
rect -276 -5851 -260 -5683
rect -348 -5867 -260 -5851
rect 245 -5683 333 -5667
rect 245 -5851 261 -5683
rect 295 -5851 333 -5683
rect 245 -5867 333 -5851
rect 1133 -5683 1221 -5667
rect 1133 -5851 1171 -5683
rect 1205 -5851 1221 -5683
rect 1133 -5867 1221 -5851
rect -1236 -5941 -1148 -5925
rect -1236 -6109 -1220 -5941
rect -1186 -6109 -1148 -5941
rect -1236 -6125 -1148 -6109
rect -348 -5941 -260 -5925
rect -348 -6109 -310 -5941
rect -276 -6109 -260 -5941
rect -348 -6125 -260 -6109
rect 245 -5941 333 -5925
rect 245 -6109 261 -5941
rect 295 -6109 333 -5941
rect 245 -6125 333 -6109
rect 1133 -5941 1221 -5925
rect 1133 -6109 1171 -5941
rect 1205 -6109 1221 -5941
rect 1133 -6125 1221 -6109
rect -1236 -6199 -1148 -6183
rect -1236 -6367 -1220 -6199
rect -1186 -6367 -1148 -6199
rect -1236 -6383 -1148 -6367
rect -348 -6199 -260 -6183
rect -348 -6367 -310 -6199
rect -276 -6367 -260 -6199
rect -348 -6383 -260 -6367
rect 245 -6199 333 -6183
rect 245 -6367 261 -6199
rect 295 -6367 333 -6199
rect 245 -6383 333 -6367
rect 1133 -6199 1221 -6183
rect 1133 -6367 1171 -6199
rect 1205 -6367 1221 -6199
rect 1133 -6383 1221 -6367
rect -1236 -6457 -1148 -6441
rect -1236 -6625 -1220 -6457
rect -1186 -6625 -1148 -6457
rect -1236 -6641 -1148 -6625
rect -348 -6457 -260 -6441
rect -348 -6625 -310 -6457
rect -276 -6625 -260 -6457
rect -348 -6641 -260 -6625
rect 245 -6457 333 -6441
rect 245 -6625 261 -6457
rect 295 -6625 333 -6457
rect 245 -6641 333 -6625
rect 1133 -6457 1221 -6441
rect 1133 -6625 1171 -6457
rect 1205 -6625 1221 -6457
rect 1133 -6641 1221 -6625
rect -1236 -6715 -1148 -6699
rect -1236 -6883 -1220 -6715
rect -1186 -6883 -1148 -6715
rect -1236 -6899 -1148 -6883
rect -348 -6715 -260 -6699
rect -348 -6883 -310 -6715
rect -276 -6883 -260 -6715
rect -348 -6899 -260 -6883
rect 245 -6715 333 -6699
rect 245 -6883 261 -6715
rect 295 -6883 333 -6715
rect 245 -6899 333 -6883
rect 1133 -6715 1221 -6699
rect 1133 -6883 1171 -6715
rect 1205 -6883 1221 -6715
rect 1133 -6899 1221 -6883
rect -1236 -6973 -1148 -6957
rect -1236 -7141 -1220 -6973
rect -1186 -7141 -1148 -6973
rect -1236 -7157 -1148 -7141
rect -348 -6973 -260 -6957
rect -348 -7141 -310 -6973
rect -276 -7141 -260 -6973
rect -348 -7157 -260 -7141
rect 245 -6973 333 -6957
rect 245 -7141 261 -6973
rect 295 -7141 333 -6973
rect 245 -7157 333 -7141
rect 1133 -6973 1221 -6957
rect 1133 -7141 1171 -6973
rect 1205 -7141 1221 -6973
rect 1133 -7157 1221 -7141
rect -1236 -7231 -1148 -7215
rect -1236 -7399 -1220 -7231
rect -1186 -7399 -1148 -7231
rect -1236 -7415 -1148 -7399
rect -348 -7231 -260 -7215
rect -348 -7399 -310 -7231
rect -276 -7399 -260 -7231
rect -348 -7415 -260 -7399
rect 245 -7231 333 -7215
rect 245 -7399 261 -7231
rect 295 -7399 333 -7231
rect 245 -7415 333 -7399
rect 1133 -7231 1221 -7215
rect 1133 -7399 1171 -7231
rect 1205 -7399 1221 -7231
rect 1133 -7415 1221 -7399
rect -1236 -7489 -1148 -7473
rect -1236 -7657 -1220 -7489
rect -1186 -7657 -1148 -7489
rect -1236 -7673 -1148 -7657
rect -348 -7489 -260 -7473
rect -348 -7657 -310 -7489
rect -276 -7657 -260 -7489
rect -348 -7673 -260 -7657
rect 245 -7489 333 -7473
rect 245 -7657 261 -7489
rect 295 -7657 333 -7489
rect 245 -7673 333 -7657
rect 1133 -7489 1221 -7473
rect 1133 -7657 1171 -7489
rect 1205 -7657 1221 -7489
rect 1133 -7673 1221 -7657
rect -1236 -7747 -1148 -7731
rect -1236 -7915 -1220 -7747
rect -1186 -7915 -1148 -7747
rect -1236 -7931 -1148 -7915
rect -348 -7747 -260 -7731
rect -348 -7915 -310 -7747
rect -276 -7915 -260 -7747
rect -348 -7931 -260 -7915
rect 245 -7747 333 -7731
rect 245 -7915 261 -7747
rect 295 -7915 333 -7747
rect 245 -7931 333 -7915
rect 1133 -7747 1221 -7731
rect 1133 -7915 1171 -7747
rect 1205 -7915 1221 -7747
rect 1133 -7931 1221 -7915
rect -1236 -8005 -1148 -7989
rect -1236 -8173 -1220 -8005
rect -1186 -8173 -1148 -8005
rect -1236 -8189 -1148 -8173
rect -348 -8005 -260 -7989
rect -348 -8173 -310 -8005
rect -276 -8173 -260 -8005
rect -348 -8189 -260 -8173
rect 245 -8005 333 -7989
rect 245 -8173 261 -8005
rect 295 -8173 333 -8005
rect 245 -8189 333 -8173
rect 1133 -8005 1221 -7989
rect 1133 -8173 1171 -8005
rect 1205 -8173 1221 -8005
rect 1133 -8189 1221 -8173
rect -1236 -8263 -1148 -8247
rect -1236 -8431 -1220 -8263
rect -1186 -8431 -1148 -8263
rect -1236 -8447 -1148 -8431
rect -348 -8263 -260 -8247
rect -348 -8431 -310 -8263
rect -276 -8431 -260 -8263
rect -348 -8447 -260 -8431
rect 245 -8263 333 -8247
rect 245 -8431 261 -8263
rect 295 -8431 333 -8263
rect 245 -8447 333 -8431
rect 1133 -8263 1221 -8247
rect 1133 -8431 1171 -8263
rect 1205 -8431 1221 -8263
rect 1133 -8447 1221 -8431
rect -1236 -8521 -1148 -8505
rect -1236 -8689 -1220 -8521
rect -1186 -8689 -1148 -8521
rect -1236 -8705 -1148 -8689
rect -348 -8521 -260 -8505
rect -348 -8689 -310 -8521
rect -276 -8689 -260 -8521
rect -348 -8705 -260 -8689
rect 245 -8521 333 -8505
rect 245 -8689 261 -8521
rect 295 -8689 333 -8521
rect 245 -8705 333 -8689
rect 1133 -8521 1221 -8505
rect 1133 -8689 1171 -8521
rect 1205 -8689 1221 -8521
rect 1133 -8705 1221 -8689
rect -1236 -8779 -1148 -8763
rect -1236 -8947 -1220 -8779
rect -1186 -8947 -1148 -8779
rect -1236 -8963 -1148 -8947
rect -348 -8779 -260 -8763
rect -348 -8947 -310 -8779
rect -276 -8947 -260 -8779
rect -348 -8963 -260 -8947
rect 245 -8779 333 -8763
rect 245 -8947 261 -8779
rect 295 -8947 333 -8779
rect 245 -8963 333 -8947
rect 1133 -8779 1221 -8763
rect 1133 -8947 1171 -8779
rect 1205 -8947 1221 -8779
rect 1133 -8963 1221 -8947
rect -1236 -9037 -1148 -9021
rect -1236 -9205 -1220 -9037
rect -1186 -9205 -1148 -9037
rect -1236 -9221 -1148 -9205
rect -348 -9037 -260 -9021
rect -348 -9205 -310 -9037
rect -276 -9205 -260 -9037
rect -348 -9221 -260 -9205
rect 245 -9037 333 -9021
rect 245 -9205 261 -9037
rect 295 -9205 333 -9037
rect 245 -9221 333 -9205
rect 1133 -9037 1221 -9021
rect 1133 -9205 1171 -9037
rect 1205 -9205 1221 -9037
rect 1133 -9221 1221 -9205
rect -1236 -9295 -1148 -9279
rect -1236 -9463 -1220 -9295
rect -1186 -9463 -1148 -9295
rect -1236 -9479 -1148 -9463
rect -348 -9295 -260 -9279
rect -348 -9463 -310 -9295
rect -276 -9463 -260 -9295
rect -348 -9479 -260 -9463
rect 245 -9295 333 -9279
rect 245 -9463 261 -9295
rect 295 -9463 333 -9295
rect 245 -9479 333 -9463
rect 1133 -9295 1221 -9279
rect 1133 -9463 1171 -9295
rect 1205 -9463 1221 -9295
rect 1133 -9479 1221 -9463
rect -1236 -9553 -1148 -9537
rect -1236 -9721 -1220 -9553
rect -1186 -9721 -1148 -9553
rect -1236 -9737 -1148 -9721
rect -348 -9553 -260 -9537
rect -348 -9721 -310 -9553
rect -276 -9721 -260 -9553
rect -348 -9737 -260 -9721
rect 245 -9553 333 -9537
rect 245 -9721 261 -9553
rect 295 -9721 333 -9553
rect 245 -9737 333 -9721
rect 1133 -9553 1221 -9537
rect 1133 -9721 1171 -9553
rect 1205 -9721 1221 -9553
rect 1133 -9737 1221 -9721
rect -1236 -9811 -1148 -9795
rect -1236 -9979 -1220 -9811
rect -1186 -9979 -1148 -9811
rect -1236 -9995 -1148 -9979
rect -348 -9811 -260 -9795
rect -348 -9979 -310 -9811
rect -276 -9979 -260 -9811
rect -348 -9995 -260 -9979
rect 245 -9811 333 -9795
rect 245 -9979 261 -9811
rect 295 -9979 333 -9811
rect 245 -9995 333 -9979
rect 1133 -9811 1221 -9795
rect 1133 -9979 1171 -9811
rect 1205 -9979 1221 -9811
rect 1133 -9995 1221 -9979
rect 2382 -3072 2470 -3056
rect 2382 -3240 2398 -3072
rect 2432 -3240 2470 -3072
rect 2382 -3256 2470 -3240
rect 2670 -3072 2758 -3056
rect 2670 -3240 2708 -3072
rect 2742 -3240 2758 -3072
rect 2670 -3256 2758 -3240
rect 2382 -3330 2470 -3314
rect 2382 -3498 2398 -3330
rect 2432 -3498 2470 -3330
rect 2382 -3514 2470 -3498
rect 2670 -3330 2758 -3314
rect 2670 -3498 2708 -3330
rect 2742 -3498 2758 -3330
rect 2670 -3514 2758 -3498
rect 2382 -3588 2470 -3572
rect 2382 -3756 2398 -3588
rect 2432 -3756 2470 -3588
rect 2382 -3772 2470 -3756
rect 2670 -3588 2758 -3572
rect 2670 -3756 2708 -3588
rect 2742 -3756 2758 -3588
rect 2670 -3772 2758 -3756
rect 2382 -3846 2470 -3830
rect 2382 -4014 2398 -3846
rect 2432 -4014 2470 -3846
rect 2382 -4030 2470 -4014
rect 2670 -3846 2758 -3830
rect 2670 -4014 2708 -3846
rect 2742 -4014 2758 -3846
rect 2670 -4030 2758 -4014
rect 2382 -4104 2470 -4088
rect 2382 -4272 2398 -4104
rect 2432 -4272 2470 -4104
rect 2382 -4288 2470 -4272
rect 2670 -4104 2758 -4088
rect 2670 -4272 2708 -4104
rect 2742 -4272 2758 -4104
rect 2670 -4288 2758 -4272
rect 2382 -4362 2470 -4346
rect 2382 -4530 2398 -4362
rect 2432 -4530 2470 -4362
rect 2382 -4546 2470 -4530
rect 2670 -4362 2758 -4346
rect 2670 -4530 2708 -4362
rect 2742 -4530 2758 -4362
rect 2670 -4546 2758 -4530
rect 2382 -4620 2470 -4604
rect 2382 -4788 2398 -4620
rect 2432 -4788 2470 -4620
rect 2382 -4804 2470 -4788
rect 2670 -4620 2758 -4604
rect 2670 -4788 2708 -4620
rect 2742 -4788 2758 -4620
rect 2670 -4804 2758 -4788
rect 2382 -4878 2470 -4862
rect 2382 -5046 2398 -4878
rect 2432 -5046 2470 -4878
rect 2382 -5062 2470 -5046
rect 2670 -4878 2758 -4862
rect 2670 -5046 2708 -4878
rect 2742 -5046 2758 -4878
rect 2670 -5062 2758 -5046
rect 2382 -5136 2470 -5120
rect 2382 -5304 2398 -5136
rect 2432 -5304 2470 -5136
rect 2382 -5320 2470 -5304
rect 2670 -5136 2758 -5120
rect 2670 -5304 2708 -5136
rect 2742 -5304 2758 -5136
rect 2670 -5320 2758 -5304
rect 2382 -5394 2470 -5378
rect 2382 -5562 2398 -5394
rect 2432 -5562 2470 -5394
rect 2382 -5578 2470 -5562
rect 2670 -5394 2758 -5378
rect 2670 -5562 2708 -5394
rect 2742 -5562 2758 -5394
rect 2670 -5578 2758 -5562
rect 2382 -5652 2470 -5636
rect 2382 -5820 2398 -5652
rect 2432 -5820 2470 -5652
rect 2382 -5836 2470 -5820
rect 2670 -5652 2758 -5636
rect 2670 -5820 2708 -5652
rect 2742 -5820 2758 -5652
rect 2670 -5836 2758 -5820
rect 2382 -5910 2470 -5894
rect 2382 -6078 2398 -5910
rect 2432 -6078 2470 -5910
rect 2382 -6094 2470 -6078
rect 2670 -5910 2758 -5894
rect 2670 -6078 2708 -5910
rect 2742 -6078 2758 -5910
rect 2670 -6094 2758 -6078
rect 2382 -6168 2470 -6152
rect 2382 -6336 2398 -6168
rect 2432 -6336 2470 -6168
rect 2382 -6352 2470 -6336
rect 2670 -6168 2758 -6152
rect 2670 -6336 2708 -6168
rect 2742 -6336 2758 -6168
rect 2670 -6352 2758 -6336
rect 2382 -6426 2470 -6410
rect 2382 -6594 2398 -6426
rect 2432 -6594 2470 -6426
rect 2382 -6610 2470 -6594
rect 2670 -6426 2758 -6410
rect 2670 -6594 2708 -6426
rect 2742 -6594 2758 -6426
rect 2670 -6610 2758 -6594
rect 2382 -6684 2470 -6668
rect 2382 -6852 2398 -6684
rect 2432 -6852 2470 -6684
rect 2382 -6868 2470 -6852
rect 2670 -6684 2758 -6668
rect 2670 -6852 2708 -6684
rect 2742 -6852 2758 -6684
rect 2670 -6868 2758 -6852
rect 2382 -6942 2470 -6926
rect 2382 -7110 2398 -6942
rect 2432 -7110 2470 -6942
rect 2382 -7126 2470 -7110
rect 2670 -6942 2758 -6926
rect 2670 -7110 2708 -6942
rect 2742 -7110 2758 -6942
rect 2670 -7126 2758 -7110
rect 2382 -7200 2470 -7184
rect 2382 -7368 2398 -7200
rect 2432 -7368 2470 -7200
rect 2382 -7384 2470 -7368
rect 2670 -7200 2758 -7184
rect 2670 -7368 2708 -7200
rect 2742 -7368 2758 -7200
rect 2670 -7384 2758 -7368
rect 2382 -7458 2470 -7442
rect 2382 -7626 2398 -7458
rect 2432 -7626 2470 -7458
rect 2382 -7642 2470 -7626
rect 2670 -7458 2758 -7442
rect 2670 -7626 2708 -7458
rect 2742 -7626 2758 -7458
rect 2670 -7642 2758 -7626
rect 2382 -7716 2470 -7700
rect 2382 -7884 2398 -7716
rect 2432 -7884 2470 -7716
rect 2382 -7900 2470 -7884
rect 2670 -7716 2758 -7700
rect 2670 -7884 2708 -7716
rect 2742 -7884 2758 -7716
rect 2670 -7900 2758 -7884
rect 2382 -7974 2470 -7958
rect 2382 -8142 2398 -7974
rect 2432 -8142 2470 -7974
rect 2382 -8158 2470 -8142
rect 2670 -7974 2758 -7958
rect 2670 -8142 2708 -7974
rect 2742 -8142 2758 -7974
rect 2670 -8158 2758 -8142
rect 3160 -3007 3257 -2991
rect 3160 -3375 3176 -3007
rect 3210 -3375 3257 -3007
rect 3160 -3391 3257 -3375
rect 3457 -3007 3554 -2991
rect 3457 -3375 3504 -3007
rect 3538 -3375 3554 -3007
rect 3457 -3391 3554 -3375
rect 3160 -3588 3257 -3572
rect 3160 -3956 3176 -3588
rect 3210 -3956 3257 -3588
rect 3160 -3972 3257 -3956
rect 3457 -3588 3554 -3572
rect 3457 -3956 3504 -3588
rect 3538 -3956 3554 -3588
rect 3457 -3972 3554 -3956
rect 8952 -2697 9040 -2681
rect 8952 -2965 8968 -2697
rect 9002 -2965 9040 -2697
rect 8952 -2981 9040 -2965
rect 10140 -2697 10228 -2681
rect 10140 -2965 10178 -2697
rect 10212 -2965 10228 -2697
rect 10140 -2981 10228 -2965
rect 8952 -3055 9040 -3039
rect 8952 -3323 8968 -3055
rect 9002 -3323 9040 -3055
rect 8952 -3339 9040 -3323
rect 10140 -3055 10228 -3039
rect 10140 -3323 10178 -3055
rect 10212 -3323 10228 -3055
rect 10140 -3339 10228 -3323
rect 3160 -4878 3257 -4862
rect 3160 -5246 3176 -4878
rect 3210 -5246 3257 -4878
rect 3160 -5262 3257 -5246
rect 3457 -4878 3554 -4862
rect 3457 -5246 3504 -4878
rect 3538 -5246 3554 -4878
rect 3457 -5262 3554 -5246
rect 3160 -6168 3257 -6152
rect 3160 -6536 3176 -6168
rect 3210 -6536 3257 -6168
rect 3160 -6552 3257 -6536
rect 3457 -6168 3554 -6152
rect 3457 -6536 3504 -6168
rect 3538 -6536 3554 -6168
rect 3457 -6552 3554 -6536
rect 3160 -7458 3257 -7442
rect 3160 -7826 3176 -7458
rect 3210 -7826 3257 -7458
rect 3160 -7842 3257 -7826
rect 3457 -7458 3554 -7442
rect 3457 -7826 3504 -7458
rect 3538 -7826 3554 -7458
rect 3457 -7842 3554 -7826
rect 3160 -8546 3257 -8530
rect 3160 -8714 3176 -8546
rect 3210 -8714 3257 -8546
rect 3160 -8730 3257 -8714
rect 3457 -8546 3554 -8530
rect 3457 -8714 3504 -8546
rect 3538 -8714 3554 -8546
rect 3457 -8730 3554 -8714
rect 3160 -8804 3257 -8788
rect 3160 -8972 3176 -8804
rect 3210 -8972 3257 -8804
rect 3160 -8988 3257 -8972
rect 3457 -8804 3554 -8788
rect 3457 -8972 3504 -8804
rect 3538 -8972 3554 -8804
rect 3457 -8988 3554 -8972
rect 3160 -9271 3257 -9255
rect 3160 -9639 3176 -9271
rect 3210 -9639 3257 -9271
rect 3160 -9655 3257 -9639
rect 3357 -9271 3454 -9255
rect 3357 -9639 3404 -9271
rect 3438 -9639 3454 -9271
rect 3357 -9655 3454 -9639
rect 3160 -9729 3257 -9713
rect 3160 -10097 3176 -9729
rect 3210 -10097 3257 -9729
rect 3160 -10113 3257 -10097
rect 3357 -9729 3454 -9713
rect 3357 -10097 3404 -9729
rect 3438 -10097 3454 -9729
rect 3357 -10113 3454 -10097
<< polycont >>
rect -9886 5114 -6318 5148
rect -6228 5114 -2660 5148
rect -9886 4626 -6318 4660
rect -6228 4626 -2660 4660
rect -9886 4138 -6318 4172
rect -6228 4138 -2660 4172
rect -10149 640 -10115 1608
rect -9439 640 -9405 1608
rect -8676 3233 -6308 3267
rect -6218 3233 -3850 3267
rect -8676 1923 -6308 1957
rect -6218 1923 -3850 1957
rect -8677 1358 -6309 1392
rect -6219 1358 -3851 1392
rect -8677 48 -6309 82
rect -6219 48 -3851 82
rect -1414 7190 -1066 7224
rect -976 7190 -628 7224
rect -538 7190 -190 7224
rect -100 7190 248 7224
rect -1414 4062 -1066 4096
rect -976 4062 -628 4096
rect -538 4062 -190 4096
rect -100 4062 248 4096
rect -1414 3213 -1066 3247
rect -976 3213 -628 3247
rect -538 3213 -190 3247
rect -100 3213 248 3247
rect -1414 85 -1066 119
rect -976 85 -628 119
rect -538 85 -190 119
rect -100 85 248 119
rect 3415 1659 3743 1693
rect 3833 1659 4161 1693
rect 4251 1659 4579 1693
rect 4669 1659 4997 1693
rect 3415 131 3743 165
rect 3833 131 4161 165
rect 4251 131 4579 165
rect 4669 131 4997 165
rect 7508 2204 8476 2238
rect 8566 2204 9534 2238
rect 9624 2204 10592 2238
rect 10682 2204 11650 2238
rect 7508 1576 8476 1610
rect 8566 1576 9534 1610
rect 9624 1576 10592 1610
rect 10682 1576 11650 1610
rect 7508 1042 8476 1076
rect 8566 1042 9534 1076
rect 9624 1042 10592 1076
rect 10682 1042 11650 1076
rect 7508 414 8476 448
rect 8566 414 9534 448
rect 9624 414 10592 448
rect 10682 414 11650 448
rect -1404 -822 444 -788
rect 534 -822 2382 -788
rect 2472 -822 4320 -788
rect 4410 -822 6258 -788
rect -1404 -1232 444 -1198
rect 534 -1232 2382 -1198
rect 2472 -1232 4320 -1198
rect 4410 -1232 6258 -1198
rect -1404 -1642 444 -1608
rect 534 -1642 2382 -1608
rect 2472 -1642 4320 -1608
rect 4410 -1642 6258 -1608
rect 8693 -252 9061 -218
rect 9151 -252 9519 -218
rect 9609 -252 9977 -218
rect 10067 -252 10435 -218
rect 8693 -962 9061 -928
rect 9151 -962 9519 -928
rect 9609 -962 9977 -928
rect 10067 -962 10435 -928
rect 8693 -1459 9061 -1425
rect 9151 -1459 9519 -1425
rect 9609 -1459 9977 -1425
rect 10067 -1459 10435 -1425
rect 8693 -2169 9061 -2135
rect 9151 -2169 9519 -2135
rect 9609 -2169 9977 -2135
rect 10067 -2169 10435 -2135
rect 11841 -361 11879 -327
rect 11841 -1009 11879 -975
rect 12197 -361 12235 -327
rect 12197 -1009 12235 -975
rect 11863 -1375 11897 -1341
rect 12219 -1375 12253 -1341
rect 11863 -1685 11897 -1651
rect 12219 -1685 12253 -1651
rect -1220 -4045 -1186 -3877
rect -310 -4045 -276 -3877
rect 261 -4045 295 -3877
rect 1171 -4045 1205 -3877
rect -1220 -4303 -1186 -4135
rect -310 -4303 -276 -4135
rect 261 -4303 295 -4135
rect 1171 -4303 1205 -4135
rect -1220 -4561 -1186 -4393
rect -310 -4561 -276 -4393
rect 261 -4561 295 -4393
rect 1171 -4561 1205 -4393
rect -1220 -4819 -1186 -4651
rect -310 -4819 -276 -4651
rect 261 -4819 295 -4651
rect 1171 -4819 1205 -4651
rect -1220 -5077 -1186 -4909
rect -310 -5077 -276 -4909
rect 261 -5077 295 -4909
rect 1171 -5077 1205 -4909
rect -1220 -5335 -1186 -5167
rect -310 -5335 -276 -5167
rect 261 -5335 295 -5167
rect 1171 -5335 1205 -5167
rect -1220 -5593 -1186 -5425
rect -310 -5593 -276 -5425
rect 261 -5593 295 -5425
rect 1171 -5593 1205 -5425
rect -1220 -5851 -1186 -5683
rect -310 -5851 -276 -5683
rect 261 -5851 295 -5683
rect 1171 -5851 1205 -5683
rect -1220 -6109 -1186 -5941
rect -310 -6109 -276 -5941
rect 261 -6109 295 -5941
rect 1171 -6109 1205 -5941
rect -1220 -6367 -1186 -6199
rect -310 -6367 -276 -6199
rect 261 -6367 295 -6199
rect 1171 -6367 1205 -6199
rect -1220 -6625 -1186 -6457
rect -310 -6625 -276 -6457
rect 261 -6625 295 -6457
rect 1171 -6625 1205 -6457
rect -1220 -6883 -1186 -6715
rect -310 -6883 -276 -6715
rect 261 -6883 295 -6715
rect 1171 -6883 1205 -6715
rect -1220 -7141 -1186 -6973
rect -310 -7141 -276 -6973
rect 261 -7141 295 -6973
rect 1171 -7141 1205 -6973
rect -1220 -7399 -1186 -7231
rect -310 -7399 -276 -7231
rect 261 -7399 295 -7231
rect 1171 -7399 1205 -7231
rect -1220 -7657 -1186 -7489
rect -310 -7657 -276 -7489
rect 261 -7657 295 -7489
rect 1171 -7657 1205 -7489
rect -1220 -7915 -1186 -7747
rect -310 -7915 -276 -7747
rect 261 -7915 295 -7747
rect 1171 -7915 1205 -7747
rect -1220 -8173 -1186 -8005
rect -310 -8173 -276 -8005
rect 261 -8173 295 -8005
rect 1171 -8173 1205 -8005
rect -1220 -8431 -1186 -8263
rect -310 -8431 -276 -8263
rect 261 -8431 295 -8263
rect 1171 -8431 1205 -8263
rect -1220 -8689 -1186 -8521
rect -310 -8689 -276 -8521
rect 261 -8689 295 -8521
rect 1171 -8689 1205 -8521
rect -1220 -8947 -1186 -8779
rect -310 -8947 -276 -8779
rect 261 -8947 295 -8779
rect 1171 -8947 1205 -8779
rect -1220 -9205 -1186 -9037
rect -310 -9205 -276 -9037
rect 261 -9205 295 -9037
rect 1171 -9205 1205 -9037
rect -1220 -9463 -1186 -9295
rect -310 -9463 -276 -9295
rect 261 -9463 295 -9295
rect 1171 -9463 1205 -9295
rect -1220 -9721 -1186 -9553
rect -310 -9721 -276 -9553
rect 261 -9721 295 -9553
rect 1171 -9721 1205 -9553
rect -1220 -9979 -1186 -9811
rect -310 -9979 -276 -9811
rect 261 -9979 295 -9811
rect 1171 -9979 1205 -9811
rect 2398 -3240 2432 -3072
rect 2708 -3240 2742 -3072
rect 2398 -3498 2432 -3330
rect 2708 -3498 2742 -3330
rect 2398 -3756 2432 -3588
rect 2708 -3756 2742 -3588
rect 2398 -4014 2432 -3846
rect 2708 -4014 2742 -3846
rect 2398 -4272 2432 -4104
rect 2708 -4272 2742 -4104
rect 2398 -4530 2432 -4362
rect 2708 -4530 2742 -4362
rect 2398 -4788 2432 -4620
rect 2708 -4788 2742 -4620
rect 2398 -5046 2432 -4878
rect 2708 -5046 2742 -4878
rect 2398 -5304 2432 -5136
rect 2708 -5304 2742 -5136
rect 2398 -5562 2432 -5394
rect 2708 -5562 2742 -5394
rect 2398 -5820 2432 -5652
rect 2708 -5820 2742 -5652
rect 2398 -6078 2432 -5910
rect 2708 -6078 2742 -5910
rect 2398 -6336 2432 -6168
rect 2708 -6336 2742 -6168
rect 2398 -6594 2432 -6426
rect 2708 -6594 2742 -6426
rect 2398 -6852 2432 -6684
rect 2708 -6852 2742 -6684
rect 2398 -7110 2432 -6942
rect 2708 -7110 2742 -6942
rect 2398 -7368 2432 -7200
rect 2708 -7368 2742 -7200
rect 2398 -7626 2432 -7458
rect 2708 -7626 2742 -7458
rect 2398 -7884 2432 -7716
rect 2708 -7884 2742 -7716
rect 2398 -8142 2432 -7974
rect 2708 -8142 2742 -7974
rect 3176 -3375 3210 -3007
rect 3504 -3375 3538 -3007
rect 3176 -3956 3210 -3588
rect 3504 -3956 3538 -3588
rect 8968 -2965 9002 -2697
rect 10178 -2965 10212 -2697
rect 8968 -3323 9002 -3055
rect 10178 -3323 10212 -3055
rect 3176 -5246 3210 -4878
rect 3504 -5246 3538 -4878
rect 3176 -6536 3210 -6168
rect 3504 -6536 3538 -6168
rect 3176 -7826 3210 -7458
rect 3504 -7826 3538 -7458
rect 3176 -8714 3210 -8546
rect 3504 -8714 3538 -8546
rect 3176 -8972 3210 -8804
rect 3504 -8972 3538 -8804
rect 3176 -9639 3210 -9271
rect 3404 -9639 3438 -9271
rect 3176 -10097 3210 -9729
rect 3404 -10097 3438 -9729
<< xpolycontact >>
rect 11275 -2439 11707 -2369
rect 11915 -2439 12347 -2369
<< xpolyres >>
rect 11707 -2439 11915 -2369
<< locali >>
rect -1848 7627 817 7640
rect -10397 5505 -2221 5541
rect -10397 5416 -10213 5505
rect -2415 5416 -2221 5505
rect -10397 5360 -2221 5416
rect -10397 5326 -10145 5360
rect -2457 5326 -2221 5360
rect -10397 5300 -2221 5326
rect -10397 4044 -10205 5300
rect -10171 5203 -2431 5300
rect -10171 4044 -10143 5203
rect -9902 5114 -9886 5148
rect -6318 5114 -6302 5148
rect -6244 5114 -6228 5148
rect -2660 5114 -2644 5148
rect -9948 5055 -9914 5071
rect -9948 4703 -9914 4719
rect -6290 5055 -6256 5071
rect -6290 4703 -6256 4719
rect -2632 5055 -2598 5071
rect -2632 4703 -2598 4719
rect -9902 4626 -9886 4660
rect -6318 4626 -6302 4660
rect -6244 4626 -6228 4660
rect -2660 4626 -2644 4660
rect -9948 4567 -9914 4583
rect -9948 4215 -9914 4231
rect -6290 4567 -6256 4583
rect -6290 4215 -6256 4231
rect -2632 4567 -2598 4583
rect -2632 4215 -2598 4231
rect -9902 4138 -9886 4172
rect -6318 4138 -6302 4172
rect -6244 4138 -6228 4172
rect -2660 4138 -2644 4172
rect -10397 4034 -10143 4044
rect -2397 5203 -2221 5300
rect -2397 4044 -2222 5203
rect -2431 4034 -2222 4044
rect -10397 4018 -2222 4034
rect -10397 3984 -10145 4018
rect -2457 3984 -2222 4018
rect -10397 3901 -2222 3984
rect -1848 4016 -1814 7627
rect 778 7424 817 7627
rect -1649 7406 626 7424
rect -1649 4016 -1614 7406
rect -1430 7190 -1414 7224
rect -1066 7190 -1050 7224
rect -992 7190 -976 7224
rect -628 7190 -612 7224
rect -554 7190 -538 7224
rect -190 7190 -174 7224
rect -116 7190 -100 7224
rect 248 7190 264 7224
rect -1476 7131 -1442 7147
rect -1476 4139 -1442 4155
rect -1038 7131 -1004 7147
rect -1038 4139 -1004 4155
rect -600 7131 -566 7147
rect -600 4139 -566 4155
rect -162 7131 -128 7147
rect -162 4139 -128 4155
rect 276 7131 310 7147
rect 276 4139 310 4155
rect 501 6845 626 7406
rect 660 6845 817 7424
rect 501 4365 566 6845
rect 708 4365 817 6845
rect -1430 4062 -1414 4096
rect -1066 4062 -1050 4096
rect -992 4062 -976 4096
rect -628 4062 -612 4096
rect -554 4062 -538 4096
rect -190 4062 -174 4096
rect -116 4062 -100 4096
rect 248 4062 264 4096
rect -10396 3399 -3247 3466
rect -10396 3365 -8914 3399
rect -3613 3365 -3247 3399
rect -10396 3339 -3247 3365
rect -10396 1785 -8974 3339
rect -10397 1784 -8974 1785
rect -10397 1750 -10155 1784
rect -9399 1750 -8974 1784
rect -10397 1748 -8974 1750
rect -10397 1688 -10186 1748
rect -10397 560 -10251 1688
rect -10217 560 -10186 1688
rect -9345 1688 -8974 1748
rect -10081 1636 -10065 1670
rect -9489 1636 -9473 1670
rect -10149 1608 -10115 1624
rect -10149 624 -10115 640
rect -9439 1608 -9405 1624
rect -9439 624 -9405 640
rect -10397 502 -10186 560
rect -10081 578 -10065 612
rect -9489 578 -9473 612
rect -10081 502 -9473 578
rect -9345 560 -9337 1688
rect -9303 560 -8974 1688
rect -9345 502 -8974 560
rect -10397 498 -8974 502
rect -10397 464 -10155 498
rect -9399 464 -8974 498
rect -10397 272 -8974 464
rect -10399 68 -8974 272
rect -10399 -26 -10291 68
rect -9738 -3 -8974 68
rect -8940 3326 -3587 3339
rect -8940 -3 -8920 3326
rect -8692 3233 -8676 3267
rect -6308 3233 -6292 3267
rect -6234 3233 -6218 3267
rect -3850 3233 -3834 3267
rect -8738 3183 -8704 3199
rect -8738 1991 -8704 2007
rect -6280 3183 -6246 3199
rect -6280 1991 -6246 2007
rect -3822 3183 -3788 3199
rect -3822 1991 -3788 2007
rect -8692 1923 -8676 1957
rect -6308 1923 -6292 1957
rect -6234 1923 -6218 1957
rect -3850 1923 -3834 1957
rect -8693 1358 -8677 1392
rect -6309 1358 -6293 1392
rect -6235 1358 -6219 1392
rect -3851 1358 -3835 1392
rect -8739 1308 -8705 1324
rect -8739 116 -8705 132
rect -6281 1308 -6247 1324
rect -6281 116 -6247 132
rect -3823 1308 -3789 1324
rect -3823 116 -3789 132
rect -8693 48 -8677 82
rect -6309 48 -6293 82
rect -6235 48 -6219 82
rect -3851 48 -3835 82
rect -9738 -8 -8920 -3
rect -3597 -3 -3587 3326
rect -3553 -3 -3247 3339
rect -3597 -8 -3247 -3
rect -9738 -26 -3247 -8
rect -10399 -29 -3247 -26
rect -10399 -63 -8914 -29
rect -3613 -63 -3247 -29
rect -10399 -167 -3247 -63
rect -1848 3198 -1740 4016
rect -1706 3198 -1614 4016
rect -1430 3213 -1414 3247
rect -1066 3213 -1050 3247
rect -992 3213 -976 3247
rect -628 3213 -612 3247
rect -554 3213 -538 3247
rect -190 3213 -174 3247
rect -116 3213 -100 3247
rect 248 3213 264 3247
rect -1848 22 -1797 3198
rect -1848 -154 -1798 22
rect -1649 3 -1614 3198
rect -1476 3154 -1442 3170
rect -1476 162 -1442 178
rect -1038 3154 -1004 3170
rect -1038 162 -1004 178
rect -600 3154 -566 3170
rect -600 162 -566 178
rect -162 3154 -128 3170
rect -162 162 -128 178
rect 276 3154 310 3170
rect 276 162 310 178
rect 501 2612 626 4365
rect 660 2612 817 4365
rect 501 132 582 2612
rect 724 2201 817 2612
rect 6936 2773 12066 3145
rect 6936 2772 11789 2773
rect 6936 2407 7086 2772
rect 12048 2441 12066 2773
rect 6936 2295 7148 2407
rect 724 2114 5557 2201
rect 5514 2113 5557 2114
rect 724 1735 2986 1822
rect 724 132 817 1735
rect -1430 85 -1414 119
rect -1066 85 -1050 119
rect -992 85 -976 119
rect -628 85 -612 119
rect -554 85 -538 119
rect -190 85 -174 119
rect -116 85 -100 119
rect 248 85 264 119
rect 501 3 626 132
rect -1649 -11 626 3
rect 660 -11 817 132
rect 767 -135 817 -11
rect -1848 -155 -1685 -154
rect 767 -155 803 -135
rect -1848 -162 803 -155
rect -10399 -256 -10289 -167
rect -3355 -256 -3247 -167
rect 2941 -168 2986 1735
rect 3219 1795 5237 1822
rect 3219 1761 3335 1795
rect 5077 1761 5237 1795
rect 3219 1735 5237 1761
rect 3219 1699 3283 1735
rect 3219 125 3239 1699
rect 3273 125 3283 1699
rect 5123 1699 5237 1735
rect 3399 1659 3415 1693
rect 3743 1659 3759 1693
rect 3817 1659 3833 1693
rect 4161 1659 4177 1693
rect 4235 1659 4251 1693
rect 4579 1659 4595 1693
rect 4653 1659 4669 1693
rect 4997 1659 5013 1693
rect 3353 1600 3387 1616
rect 3353 208 3387 224
rect 3771 1600 3805 1616
rect 3771 208 3805 224
rect 4189 1600 4223 1616
rect 4189 208 4223 224
rect 4607 1600 4641 1616
rect 4607 208 4641 224
rect 5025 1600 5059 1616
rect 5025 208 5059 224
rect 3399 131 3415 165
rect 3743 131 3759 165
rect 3817 131 3833 165
rect 4161 131 4177 165
rect 4235 131 4251 165
rect 4579 131 4595 165
rect 4653 131 4669 165
rect 4997 131 5013 165
rect 3219 92 3283 125
rect 5123 125 5139 1699
rect 5173 306 5237 1699
rect 5524 306 5557 2113
rect 5173 125 5557 306
rect 5123 92 5557 125
rect 3219 72 5557 92
rect 7127 115 7148 2295
rect 11890 2407 11932 2408
rect 7265 2295 11932 2407
rect 7265 239 7307 2295
rect 7492 2204 7508 2238
rect 8476 2204 8492 2238
rect 8550 2204 8566 2238
rect 9534 2204 9550 2238
rect 9608 2204 9624 2238
rect 10592 2204 10608 2238
rect 10666 2204 10682 2238
rect 11650 2204 11666 2238
rect 7446 2145 7480 2161
rect 7446 1653 7480 1669
rect 8504 2145 8538 2161
rect 8504 1653 8538 1669
rect 9562 2145 9596 2161
rect 9562 1653 9596 1669
rect 10620 2145 10654 2161
rect 10620 1653 10654 1669
rect 11678 2145 11712 2161
rect 11678 1653 11712 1669
rect 7492 1576 7508 1610
rect 8476 1576 8492 1610
rect 8550 1576 8566 1610
rect 9534 1576 9550 1610
rect 9608 1576 9624 1610
rect 10592 1576 10608 1610
rect 10666 1576 10682 1610
rect 11650 1576 11666 1610
rect 11911 1594 11932 2295
rect 12048 2408 12069 2441
rect 12029 1594 12069 2408
rect 7492 1042 7508 1076
rect 8476 1042 8492 1076
rect 8550 1042 8566 1076
rect 9534 1042 9550 1076
rect 9608 1042 9624 1076
rect 10592 1042 10608 1076
rect 10666 1042 10682 1076
rect 11650 1042 11666 1076
rect 7446 983 7480 999
rect 7446 491 7480 507
rect 8504 983 8538 999
rect 8504 491 8538 507
rect 9562 983 9596 999
rect 9562 491 9596 507
rect 10620 983 10654 999
rect 10620 491 10654 507
rect 11678 983 11712 999
rect 11678 491 11712 507
rect 7492 414 7508 448
rect 8476 414 8492 448
rect 8550 414 8566 448
rect 9534 414 9550 448
rect 9608 414 9624 448
rect 10592 414 10608 448
rect 10666 414 10682 448
rect 11650 414 11666 448
rect 11911 239 11953 1594
rect 7265 205 11953 239
rect 11697 200 11953 205
rect 11987 200 12069 1594
rect 11697 174 12069 200
rect 11927 163 12069 174
rect 11927 140 12456 163
rect 7127 108 7183 115
rect 7127 87 11593 108
rect 7141 81 11593 87
rect 3219 66 5561 72
rect 2941 -170 3071 -168
rect 5134 -170 5561 66
rect 8479 -25 10680 0
rect 8479 -150 8506 -25
rect 10655 -122 10680 -25
rect 2941 -184 5561 -170
rect -10399 -318 -3247 -256
rect -1752 -493 6084 -456
rect -1752 -1993 -1742 -493
rect -1595 -496 6084 -493
rect 6200 -496 6655 -456
rect 6541 -530 6655 -496
rect 6200 -556 6655 -530
rect -1595 -617 6084 -605
rect 6200 -617 6567 -556
rect -1595 -643 6567 -617
rect -1595 -1721 -1574 -643
rect -1420 -822 -1404 -788
rect 444 -822 460 -788
rect 518 -822 534 -788
rect 2382 -822 2398 -788
rect 2456 -822 2472 -788
rect 4320 -822 4336 -788
rect 4394 -822 4410 -788
rect 6258 -822 6274 -788
rect -1466 -872 -1432 -856
rect -1466 -1164 -1432 -1148
rect 472 -872 506 -856
rect 472 -1164 506 -1148
rect 2410 -872 2444 -856
rect 2410 -1164 2444 -1148
rect 4348 -872 4382 -856
rect 4348 -1164 4382 -1148
rect 6286 -872 6320 -856
rect 6286 -1164 6320 -1148
rect -1420 -1232 -1404 -1198
rect 444 -1232 460 -1198
rect 518 -1232 534 -1198
rect 2382 -1232 2398 -1198
rect 2456 -1232 2472 -1198
rect 4320 -1232 4336 -1198
rect 4394 -1232 4410 -1198
rect 6258 -1232 6274 -1198
rect -1466 -1282 -1432 -1266
rect -1466 -1574 -1432 -1558
rect 472 -1282 506 -1266
rect 472 -1574 506 -1558
rect 2410 -1282 2444 -1266
rect 2410 -1574 2444 -1558
rect 4348 -1282 4382 -1266
rect 4348 -1574 4382 -1558
rect 6286 -1282 6320 -1266
rect 6286 -1574 6320 -1558
rect -1420 -1642 -1404 -1608
rect 444 -1642 460 -1608
rect 518 -1642 534 -1608
rect 2382 -1642 2398 -1608
rect 2456 -1642 2472 -1608
rect 4320 -1642 4336 -1608
rect 4394 -1642 4410 -1608
rect 6258 -1642 6274 -1608
rect 6486 -1721 6567 -643
rect -1595 -1779 6567 -1721
rect 6601 -1779 6655 -556
rect -1595 -1795 6655 -1779
rect -1501 -1796 6655 -1795
rect 6177 -1805 6655 -1796
rect 6541 -1839 6655 -1805
rect 6177 -1993 6655 -1839
rect -1752 -2010 6655 -1993
rect -1743 -2011 6655 -2010
rect 8486 -666 8506 -150
rect 8564 -150 10579 -128
rect 8564 -666 8579 -150
rect 8677 -252 8693 -218
rect 9061 -252 9077 -218
rect 9135 -252 9151 -218
rect 9519 -252 9535 -218
rect 9593 -252 9609 -218
rect 9977 -252 9993 -218
rect 10051 -252 10067 -218
rect 10435 -252 10451 -218
rect 8486 -1702 8521 -666
rect 8555 -1702 8579 -666
rect 8631 -302 8665 -286
rect 8631 -894 8665 -878
rect 9089 -302 9123 -286
rect 9089 -894 9123 -878
rect 9547 -302 9581 -286
rect 9547 -894 9581 -878
rect 10005 -302 10039 -286
rect 10005 -894 10039 -878
rect 10463 -302 10497 -286
rect 10463 -894 10497 -878
rect 8677 -962 8693 -928
rect 9061 -962 9077 -928
rect 9135 -962 9151 -928
rect 9519 -962 9535 -928
rect 9593 -962 9609 -928
rect 9977 -962 9993 -928
rect 10051 -962 10067 -928
rect 10435 -962 10451 -928
rect 8677 -1459 8693 -1425
rect 9061 -1459 9077 -1425
rect 9135 -1459 9151 -1425
rect 9519 -1459 9535 -1425
rect 9593 -1459 9609 -1425
rect 9977 -1459 9993 -1425
rect 10051 -1459 10067 -1425
rect 10435 -1459 10451 -1425
rect 8486 -2232 8497 -1702
rect 8440 -2333 8497 -2232
rect 8571 -2232 8579 -1702
rect 8631 -1509 8665 -1493
rect 8631 -2101 8665 -2085
rect 9089 -1509 9123 -1493
rect 9089 -2101 9123 -2085
rect 9547 -1509 9581 -1493
rect 9547 -2101 9581 -2085
rect 10005 -1509 10039 -1493
rect 10005 -2101 10039 -2085
rect 10463 -1509 10497 -1493
rect 10463 -2101 10497 -2085
rect 8677 -2169 8693 -2135
rect 9061 -2169 9077 -2135
rect 9135 -2169 9151 -2135
rect 9519 -2169 9535 -2135
rect 9593 -2169 9609 -2135
rect 9977 -2169 9993 -2135
rect 10051 -2169 10067 -2135
rect 10435 -2169 10451 -2135
rect 10566 -2232 10579 -150
rect 8571 -2278 10579 -2232
rect 10655 -2231 10688 -122
rect 11572 -1051 11593 81
rect 11697 -225 12456 140
rect 11697 -259 11761 -225
rect 11959 -259 12117 -225
rect 12315 -259 12456 -225
rect 11697 -278 12456 -259
rect 11697 -321 11710 -278
rect 11699 -1015 11710 -321
rect 12021 -321 12055 -278
rect 11825 -361 11841 -327
rect 11879 -361 11895 -327
rect 11779 -420 11813 -404
rect 11779 -932 11813 -916
rect 11907 -420 11941 -404
rect 11907 -932 11941 -916
rect 11825 -1009 11841 -975
rect 11879 -1009 11895 -975
rect 11697 -1051 11710 -1015
rect 11572 -1077 11710 -1051
rect 12373 -321 12456 -278
rect 12181 -361 12197 -327
rect 12235 -361 12251 -327
rect 12135 -420 12169 -404
rect 12135 -932 12169 -916
rect 12263 -420 12297 -404
rect 12263 -932 12297 -916
rect 12181 -1009 12197 -975
rect 12235 -1009 12251 -975
rect 12021 -1077 12055 -1015
rect 12373 -1015 12377 -321
rect 12411 -1015 12456 -321
rect 12373 -1077 12456 -1015
rect 11572 -1111 11761 -1077
rect 11959 -1111 12117 -1077
rect 12315 -1111 12456 -1077
rect 11572 -1134 11710 -1111
rect 12373 -1120 12456 -1111
rect 10974 -1239 12508 -1219
rect 10974 -1273 11757 -1239
rect 12356 -1273 12508 -1239
rect 10974 -1297 12508 -1273
rect 10974 -1299 11749 -1297
rect 10974 -1739 11697 -1299
rect 11731 -1739 11749 -1299
rect 12362 -1299 12508 -1297
rect 11847 -1375 11863 -1341
rect 11897 -1375 11913 -1341
rect 12203 -1375 12219 -1341
rect 12253 -1375 12269 -1341
rect 11819 -1425 11853 -1409
rect 11819 -1617 11853 -1601
rect 11907 -1425 11941 -1409
rect 11907 -1617 11941 -1601
rect 12175 -1425 12209 -1409
rect 12175 -1617 12209 -1601
rect 12263 -1425 12297 -1409
rect 12263 -1617 12297 -1601
rect 11847 -1685 11863 -1651
rect 11897 -1685 11913 -1651
rect 12203 -1685 12219 -1651
rect 12253 -1685 12269 -1651
rect 10974 -1748 11749 -1739
rect 12362 -1739 12382 -1299
rect 12416 -1739 12508 -1299
rect 12362 -1748 12508 -1739
rect 10974 -1765 12508 -1748
rect 10974 -1799 11757 -1765
rect 12356 -1799 12508 -1765
rect 10974 -1885 12508 -1799
rect 10974 -2231 10997 -1885
rect 12375 -2157 12508 -1885
rect 8571 -2312 8581 -2278
rect 10563 -2312 10579 -2278
rect 8571 -2333 10579 -2312
rect 10655 -2333 10997 -2231
rect 11117 -2239 12508 -2157
rect 11117 -2273 11241 -2239
rect 12381 -2273 12508 -2239
rect 11117 -2295 12508 -2273
rect 8440 -2570 8452 -2333
rect 11117 -2335 11179 -2295
rect 11117 -2473 11145 -2335
rect 12437 -2335 12508 -2295
rect 11117 -2503 11179 -2473
rect 3058 -2787 3602 -2786
rect 2094 -2843 2984 -2796
rect 2094 -2877 2284 -2843
rect 2866 -2877 2984 -2843
rect 2094 -2903 2984 -2877
rect 2094 -2918 2224 -2903
rect 2258 -2918 2892 -2903
rect 2094 -3645 2122 -2918
rect 1541 -3648 2122 -3645
rect -1639 -3671 2122 -3648
rect -1639 -3685 -1364 -3671
rect -1639 -10263 -1561 -3685
rect -1387 -3705 -1364 -3685
rect 1345 -3705 2122 -3671
rect -1387 -3729 2122 -3705
rect -1387 -3731 1380 -3729
rect -1387 -3764 1371 -3731
rect -1387 -10187 -1278 -3764
rect -1152 -3849 -1136 -3815
rect -360 -3849 -344 -3815
rect 329 -3849 345 -3815
rect 1121 -3849 1137 -3815
rect -1220 -3877 -1186 -3861
rect -1220 -4061 -1186 -4045
rect -310 -3877 -276 -3861
rect -310 -4061 -276 -4045
rect 261 -3877 295 -3861
rect 261 -4061 295 -4045
rect 1171 -3877 1205 -3861
rect 1171 -4061 1205 -4045
rect -1152 -4107 -1136 -4073
rect -360 -4107 -344 -4073
rect 329 -4107 345 -4073
rect 1121 -4107 1137 -4073
rect -1220 -4135 -1186 -4119
rect -1220 -4319 -1186 -4303
rect -310 -4135 -276 -4119
rect -310 -4319 -276 -4303
rect 261 -4135 295 -4119
rect 261 -4319 295 -4303
rect 1171 -4135 1205 -4119
rect 1171 -4319 1205 -4303
rect -1152 -4365 -1136 -4331
rect -360 -4365 -344 -4331
rect 329 -4365 345 -4331
rect 1121 -4365 1137 -4331
rect -1220 -4393 -1186 -4377
rect -1220 -4577 -1186 -4561
rect -310 -4393 -276 -4377
rect -310 -4577 -276 -4561
rect 261 -4393 295 -4377
rect 261 -4577 295 -4561
rect 1171 -4393 1205 -4377
rect 1171 -4577 1205 -4561
rect -1152 -4623 -1136 -4589
rect -360 -4623 -344 -4589
rect 329 -4623 345 -4589
rect 1121 -4623 1137 -4589
rect -1220 -4651 -1186 -4635
rect -1220 -4835 -1186 -4819
rect -310 -4651 -276 -4635
rect -310 -4835 -276 -4819
rect 261 -4651 295 -4635
rect 261 -4835 295 -4819
rect 1171 -4651 1205 -4635
rect 1171 -4835 1205 -4819
rect -1152 -4881 -1136 -4847
rect -360 -4881 -344 -4847
rect 329 -4881 345 -4847
rect 1121 -4881 1137 -4847
rect -1220 -4909 -1186 -4893
rect -1220 -5093 -1186 -5077
rect -310 -4909 -276 -4893
rect -310 -5093 -276 -5077
rect 261 -4909 295 -4893
rect 261 -5093 295 -5077
rect 1171 -4909 1205 -4893
rect 1171 -5093 1205 -5077
rect -1152 -5139 -1136 -5105
rect -360 -5139 -344 -5105
rect 329 -5139 345 -5105
rect 1121 -5139 1137 -5105
rect -1220 -5167 -1186 -5151
rect -1220 -5351 -1186 -5335
rect -310 -5167 -276 -5151
rect -310 -5351 -276 -5335
rect 261 -5167 295 -5151
rect 261 -5351 295 -5335
rect 1171 -5167 1205 -5151
rect 1171 -5351 1205 -5335
rect -1152 -5397 -1136 -5363
rect -360 -5397 -344 -5363
rect 329 -5397 345 -5363
rect 1121 -5397 1137 -5363
rect -1220 -5425 -1186 -5409
rect -1220 -5609 -1186 -5593
rect -310 -5425 -276 -5409
rect -310 -5609 -276 -5593
rect 261 -5425 295 -5409
rect 261 -5609 295 -5593
rect 1171 -5425 1205 -5409
rect 1171 -5609 1205 -5593
rect -1152 -5655 -1136 -5621
rect -360 -5655 -344 -5621
rect 329 -5655 345 -5621
rect 1121 -5655 1137 -5621
rect -1220 -5683 -1186 -5667
rect -1220 -5867 -1186 -5851
rect -310 -5683 -276 -5667
rect -310 -5867 -276 -5851
rect 261 -5683 295 -5667
rect 261 -5867 295 -5851
rect 1171 -5683 1205 -5667
rect 1171 -5867 1205 -5851
rect -1152 -5913 -1136 -5879
rect -360 -5913 -344 -5879
rect 329 -5913 345 -5879
rect 1121 -5913 1137 -5879
rect -1220 -5941 -1186 -5925
rect -1220 -6125 -1186 -6109
rect -310 -5941 -276 -5925
rect -310 -6125 -276 -6109
rect 261 -5941 295 -5925
rect 261 -6125 295 -6109
rect 1171 -5941 1205 -5925
rect 1171 -6125 1205 -6109
rect -1152 -6171 -1136 -6137
rect -360 -6171 -344 -6137
rect 329 -6171 345 -6137
rect 1121 -6171 1137 -6137
rect -1220 -6199 -1186 -6183
rect -1220 -6383 -1186 -6367
rect -310 -6199 -276 -6183
rect -310 -6383 -276 -6367
rect 261 -6199 295 -6183
rect 261 -6383 295 -6367
rect 1171 -6199 1205 -6183
rect 1171 -6383 1205 -6367
rect -1152 -6429 -1136 -6395
rect -360 -6429 -344 -6395
rect 329 -6429 345 -6395
rect 1121 -6429 1137 -6395
rect -1220 -6457 -1186 -6441
rect -1220 -6641 -1186 -6625
rect -310 -6457 -276 -6441
rect -310 -6641 -276 -6625
rect 261 -6457 295 -6441
rect 261 -6641 295 -6625
rect 1171 -6457 1205 -6441
rect 1171 -6641 1205 -6625
rect -1152 -6687 -1136 -6653
rect -360 -6687 -344 -6653
rect 329 -6687 345 -6653
rect 1121 -6687 1137 -6653
rect -1220 -6715 -1186 -6699
rect -1220 -6899 -1186 -6883
rect -310 -6715 -276 -6699
rect -310 -6899 -276 -6883
rect 261 -6715 295 -6699
rect 261 -6899 295 -6883
rect 1171 -6715 1205 -6699
rect 1171 -6899 1205 -6883
rect -1152 -6945 -1136 -6911
rect -360 -6945 -344 -6911
rect 329 -6945 345 -6911
rect 1121 -6945 1137 -6911
rect -1220 -6973 -1186 -6957
rect -1220 -7157 -1186 -7141
rect -310 -6973 -276 -6957
rect -310 -7157 -276 -7141
rect 261 -6973 295 -6957
rect 261 -7157 295 -7141
rect 1171 -6973 1205 -6957
rect 1171 -7157 1205 -7141
rect -1152 -7203 -1136 -7169
rect -360 -7203 -344 -7169
rect 329 -7203 345 -7169
rect 1121 -7203 1137 -7169
rect -1220 -7231 -1186 -7215
rect -1220 -7415 -1186 -7399
rect -310 -7231 -276 -7215
rect -310 -7415 -276 -7399
rect 261 -7231 295 -7215
rect 261 -7415 295 -7399
rect 1171 -7231 1205 -7215
rect 1171 -7415 1205 -7399
rect -1152 -7461 -1136 -7427
rect -360 -7461 -344 -7427
rect 329 -7461 345 -7427
rect 1121 -7461 1137 -7427
rect -1220 -7489 -1186 -7473
rect -1220 -7673 -1186 -7657
rect -310 -7489 -276 -7473
rect -310 -7673 -276 -7657
rect 261 -7489 295 -7473
rect 261 -7673 295 -7657
rect 1171 -7489 1205 -7473
rect 1171 -7673 1205 -7657
rect -1152 -7719 -1136 -7685
rect -360 -7719 -344 -7685
rect 329 -7719 345 -7685
rect 1121 -7719 1137 -7685
rect -1220 -7747 -1186 -7731
rect -1220 -7931 -1186 -7915
rect -310 -7747 -276 -7731
rect -310 -7931 -276 -7915
rect 261 -7747 295 -7731
rect 261 -7931 295 -7915
rect 1171 -7747 1205 -7731
rect 1171 -7931 1205 -7915
rect -1152 -7977 -1136 -7943
rect -360 -7977 -344 -7943
rect 329 -7977 345 -7943
rect 1121 -7977 1137 -7943
rect -1220 -8005 -1186 -7989
rect -1220 -8189 -1186 -8173
rect -310 -8005 -276 -7989
rect -310 -8189 -276 -8173
rect 261 -8005 295 -7989
rect 261 -8189 295 -8173
rect 1171 -8005 1205 -7989
rect 1171 -8189 1205 -8173
rect -1152 -8235 -1136 -8201
rect -360 -8235 -344 -8201
rect 329 -8235 345 -8201
rect 1121 -8235 1137 -8201
rect -1220 -8263 -1186 -8247
rect -1220 -8447 -1186 -8431
rect -310 -8263 -276 -8247
rect -310 -8447 -276 -8431
rect 261 -8263 295 -8247
rect 261 -8447 295 -8431
rect 1171 -8263 1205 -8247
rect 1171 -8447 1205 -8431
rect -1152 -8493 -1136 -8459
rect -360 -8493 -344 -8459
rect 329 -8493 345 -8459
rect 1121 -8493 1137 -8459
rect -1220 -8521 -1186 -8505
rect -1220 -8705 -1186 -8689
rect -310 -8521 -276 -8505
rect -310 -8705 -276 -8689
rect 261 -8521 295 -8505
rect 261 -8705 295 -8689
rect 1171 -8521 1205 -8505
rect 1171 -8705 1205 -8689
rect -1152 -8751 -1136 -8717
rect -360 -8751 -344 -8717
rect 329 -8751 345 -8717
rect 1121 -8751 1137 -8717
rect -1220 -8779 -1186 -8763
rect -1220 -8963 -1186 -8947
rect -310 -8779 -276 -8763
rect -310 -8963 -276 -8947
rect 261 -8779 295 -8763
rect 261 -8963 295 -8947
rect 1171 -8779 1205 -8763
rect 1171 -8963 1205 -8947
rect -1152 -9009 -1136 -8975
rect -360 -9009 -344 -8975
rect 329 -9009 345 -8975
rect 1121 -9009 1137 -8975
rect -1220 -9037 -1186 -9021
rect -1220 -9221 -1186 -9205
rect -310 -9037 -276 -9021
rect -310 -9221 -276 -9205
rect 261 -9037 295 -9021
rect 261 -9221 295 -9205
rect 1171 -9037 1205 -9021
rect 1171 -9221 1205 -9205
rect -1152 -9267 -1136 -9233
rect -360 -9267 -344 -9233
rect 329 -9267 345 -9233
rect 1121 -9267 1137 -9233
rect -1220 -9295 -1186 -9279
rect -1220 -9479 -1186 -9463
rect -310 -9295 -276 -9279
rect -310 -9479 -276 -9463
rect 261 -9295 295 -9279
rect 261 -9479 295 -9463
rect 1171 -9295 1205 -9279
rect 1171 -9479 1205 -9463
rect -1152 -9525 -1136 -9491
rect -360 -9525 -344 -9491
rect 329 -9525 345 -9491
rect 1121 -9525 1137 -9491
rect -1220 -9553 -1186 -9537
rect -1220 -9737 -1186 -9721
rect -310 -9553 -276 -9537
rect -310 -9737 -276 -9721
rect 261 -9553 295 -9537
rect 261 -9737 295 -9721
rect 1171 -9553 1205 -9537
rect 1171 -9737 1205 -9721
rect -1152 -9783 -1136 -9749
rect -360 -9783 -344 -9749
rect 329 -9783 345 -9749
rect 1121 -9783 1137 -9749
rect -1220 -9811 -1186 -9795
rect -1220 -9995 -1186 -9979
rect -310 -9811 -276 -9795
rect -310 -9995 -276 -9979
rect 261 -9811 295 -9795
rect 261 -9995 295 -9979
rect 1171 -9811 1205 -9795
rect 1171 -9995 1205 -9979
rect -1152 -10041 -1136 -10007
rect -360 -10041 -344 -10007
rect 329 -10041 345 -10007
rect 1121 -10041 1137 -10007
rect 1328 -10027 1371 -3764
rect 1335 -10187 1371 -10027
rect 1492 -8325 2122 -3729
rect 2313 -2919 2892 -2918
rect 2313 -8295 2350 -2919
rect 2466 -3044 2482 -3010
rect 2658 -3044 2674 -3010
rect 2398 -3072 2432 -3056
rect 2398 -3256 2432 -3240
rect 2708 -3072 2742 -3056
rect 2708 -3256 2742 -3240
rect 2466 -3302 2482 -3268
rect 2658 -3302 2674 -3268
rect 2398 -3330 2432 -3314
rect 2398 -3514 2432 -3498
rect 2708 -3330 2742 -3314
rect 2708 -3514 2742 -3498
rect 2466 -3560 2482 -3526
rect 2658 -3560 2674 -3526
rect 2398 -3588 2432 -3572
rect 2398 -3772 2432 -3756
rect 2708 -3588 2742 -3572
rect 2708 -3772 2742 -3756
rect 2466 -3818 2482 -3784
rect 2658 -3818 2674 -3784
rect 2398 -3846 2432 -3830
rect 2398 -4030 2432 -4014
rect 2708 -3846 2742 -3830
rect 2708 -4030 2742 -4014
rect 2466 -4076 2482 -4042
rect 2658 -4076 2674 -4042
rect 2398 -4104 2432 -4088
rect 2398 -4288 2432 -4272
rect 2708 -4104 2742 -4088
rect 2708 -4288 2742 -4272
rect 2466 -4334 2482 -4300
rect 2658 -4334 2674 -4300
rect 2398 -4362 2432 -4346
rect 2398 -4546 2432 -4530
rect 2708 -4362 2742 -4346
rect 2708 -4546 2742 -4530
rect 2466 -4592 2482 -4558
rect 2658 -4592 2674 -4558
rect 2398 -4620 2432 -4604
rect 2398 -4804 2432 -4788
rect 2708 -4620 2742 -4604
rect 2708 -4804 2742 -4788
rect 2466 -4850 2482 -4816
rect 2658 -4850 2674 -4816
rect 2398 -4878 2432 -4862
rect 2398 -5062 2432 -5046
rect 2708 -4878 2742 -4862
rect 2708 -5062 2742 -5046
rect 2466 -5108 2482 -5074
rect 2658 -5108 2674 -5074
rect 2398 -5136 2432 -5120
rect 2398 -5320 2432 -5304
rect 2708 -5136 2742 -5120
rect 2708 -5320 2742 -5304
rect 2466 -5366 2482 -5332
rect 2658 -5366 2674 -5332
rect 2398 -5394 2432 -5378
rect 2398 -5578 2432 -5562
rect 2708 -5394 2742 -5378
rect 2708 -5578 2742 -5562
rect 2466 -5624 2482 -5590
rect 2658 -5624 2674 -5590
rect 2398 -5652 2432 -5636
rect 2398 -5836 2432 -5820
rect 2708 -5652 2742 -5636
rect 2708 -5836 2742 -5820
rect 2466 -5882 2482 -5848
rect 2658 -5882 2674 -5848
rect 2398 -5910 2432 -5894
rect 2398 -6094 2432 -6078
rect 2708 -5910 2742 -5894
rect 2708 -6094 2742 -6078
rect 2466 -6140 2482 -6106
rect 2658 -6140 2674 -6106
rect 2398 -6168 2432 -6152
rect 2398 -6352 2432 -6336
rect 2708 -6168 2742 -6152
rect 2708 -6352 2742 -6336
rect 2466 -6398 2482 -6364
rect 2658 -6398 2674 -6364
rect 2398 -6426 2432 -6410
rect 2398 -6610 2432 -6594
rect 2708 -6426 2742 -6410
rect 2708 -6610 2742 -6594
rect 2466 -6656 2482 -6622
rect 2658 -6656 2674 -6622
rect 2398 -6684 2432 -6668
rect 2398 -6868 2432 -6852
rect 2708 -6684 2742 -6668
rect 2708 -6868 2742 -6852
rect 2466 -6914 2482 -6880
rect 2658 -6914 2674 -6880
rect 2398 -6942 2432 -6926
rect 2398 -7126 2432 -7110
rect 2708 -6942 2742 -6926
rect 2708 -7126 2742 -7110
rect 2466 -7172 2482 -7138
rect 2658 -7172 2674 -7138
rect 2398 -7200 2432 -7184
rect 2398 -7384 2432 -7368
rect 2708 -7200 2742 -7184
rect 2708 -7384 2742 -7368
rect 2466 -7430 2482 -7396
rect 2658 -7430 2674 -7396
rect 2398 -7458 2432 -7442
rect 2398 -7642 2432 -7626
rect 2708 -7458 2742 -7442
rect 2708 -7642 2742 -7626
rect 2466 -7688 2482 -7654
rect 2658 -7688 2674 -7654
rect 2398 -7716 2432 -7700
rect 2398 -7900 2432 -7884
rect 2708 -7716 2742 -7700
rect 2708 -7900 2742 -7884
rect 2466 -7946 2482 -7912
rect 2658 -7946 2674 -7912
rect 2398 -7974 2432 -7958
rect 2398 -8158 2432 -8142
rect 2708 -7974 2742 -7958
rect 2708 -8158 2742 -8142
rect 2466 -8204 2482 -8170
rect 2658 -8204 2674 -8170
rect 2845 -8295 2892 -2919
rect 2313 -8311 2892 -8295
rect 2926 -8311 2984 -2903
rect 3058 -2835 4010 -2787
rect 3058 -2869 3158 -2835
rect 3582 -2869 4010 -2835
rect 3058 -2890 4010 -2869
rect 3058 -2895 3137 -2890
rect 3058 -4059 3098 -2895
rect 3132 -4059 3137 -2895
rect 3586 -2895 4010 -2890
rect 3253 -2979 3269 -2945
rect 3445 -2979 3461 -2945
rect 3176 -3007 3210 -2991
rect 3176 -3391 3210 -3375
rect 3504 -3007 3538 -2991
rect 3504 -3391 3538 -3375
rect 3253 -3437 3269 -3403
rect 3445 -3437 3461 -3403
rect 3253 -3560 3269 -3526
rect 3445 -3560 3461 -3526
rect 3176 -3588 3210 -3572
rect 3176 -3972 3210 -3956
rect 3504 -3588 3538 -3572
rect 3504 -3972 3538 -3956
rect 3253 -4018 3269 -3984
rect 3445 -4018 3461 -3984
rect 3058 -4073 3137 -4059
rect 3586 -4059 3608 -2895
rect 3642 -2900 4010 -2895
rect 3642 -4059 3716 -2900
rect 3586 -4073 3716 -4059
rect 3058 -4085 3716 -4073
rect 3058 -4119 3158 -4085
rect 3582 -4119 3716 -4085
rect 3058 -4156 3716 -4119
rect 3060 -4158 3716 -4156
rect 3224 -4666 3716 -4158
rect 3049 -4702 3716 -4666
rect 3049 -4736 3170 -4702
rect 3544 -4736 3716 -4702
rect 3049 -4762 3716 -4736
rect 3049 -4798 3132 -4762
rect 3585 -4763 3716 -4762
rect 3049 -5326 3074 -4798
rect 3108 -5326 3132 -4798
rect 3586 -4798 3716 -4763
rect 3253 -4850 3269 -4816
rect 3445 -4850 3461 -4816
rect 3176 -4878 3210 -4862
rect 3176 -5262 3210 -5246
rect 3504 -4878 3538 -4862
rect 3504 -5262 3538 -5246
rect 3586 -5263 3606 -4798
rect 3253 -5308 3269 -5274
rect 3445 -5308 3461 -5274
rect 3049 -5359 3132 -5326
rect 3585 -5326 3606 -5263
rect 3640 -5326 3716 -4798
rect 3585 -5359 3716 -5326
rect 3049 -5388 3716 -5359
rect 3049 -5422 3170 -5388
rect 3544 -5422 3716 -5388
rect 3049 -5450 3716 -5422
rect 3224 -5956 3716 -5450
rect 3058 -5992 3716 -5956
rect 3058 -6026 3170 -5992
rect 3544 -6026 3716 -5992
rect 3058 -6036 3716 -6026
rect 3058 -6088 3134 -6036
rect 3058 -6616 3074 -6088
rect 3108 -6616 3134 -6088
rect 3586 -6088 3716 -6036
rect 3253 -6140 3269 -6106
rect 3445 -6140 3461 -6106
rect 3176 -6168 3210 -6152
rect 3176 -6552 3210 -6536
rect 3504 -6168 3538 -6152
rect 3504 -6552 3538 -6536
rect 3253 -6598 3269 -6564
rect 3445 -6598 3461 -6564
rect 3058 -6657 3134 -6616
rect 3586 -6616 3606 -6088
rect 3640 -6616 3716 -6088
rect 3586 -6657 3716 -6616
rect 3058 -6678 3716 -6657
rect 3058 -6712 3170 -6678
rect 3544 -6712 3716 -6678
rect 3058 -6742 3716 -6712
rect 3058 -6746 3134 -6742
rect 3052 -7257 3120 -7256
rect 3236 -7257 3716 -6742
rect 3052 -7282 3716 -7257
rect 3052 -7316 3170 -7282
rect 3544 -7316 3716 -7282
rect 3052 -7335 3716 -7316
rect 3052 -7378 3120 -7335
rect 3052 -7906 3074 -7378
rect 3108 -7906 3120 -7378
rect 3586 -7378 3716 -7335
rect 3253 -7430 3269 -7396
rect 3445 -7430 3461 -7396
rect 3176 -7458 3210 -7442
rect 3176 -7842 3210 -7826
rect 3504 -7458 3538 -7442
rect 3504 -7842 3538 -7826
rect 3253 -7888 3269 -7854
rect 3445 -7888 3461 -7854
rect 3052 -7947 3120 -7906
rect 3586 -7906 3606 -7378
rect 3640 -7895 3716 -7378
rect 3855 -7895 4010 -2900
rect 8443 -3760 8452 -2570
rect 8790 -2521 10341 -2503
rect 8790 -2555 8962 -2521
rect 10218 -2555 10341 -2521
rect 8790 -2570 10341 -2555
rect 8790 -2617 8926 -2570
rect 8790 -3403 8866 -2617
rect 8900 -3403 8926 -2617
rect 10280 -2617 10341 -2570
rect 9036 -2669 9052 -2635
rect 10128 -2669 10144 -2635
rect 8968 -2697 9002 -2681
rect 8968 -2981 9002 -2965
rect 10178 -2697 10212 -2681
rect 10178 -2981 10212 -2965
rect 9036 -3027 9052 -2993
rect 10128 -3027 10144 -2993
rect 8968 -3055 9002 -3039
rect 8968 -3339 9002 -3323
rect 10178 -3055 10212 -3039
rect 10178 -3339 10212 -3323
rect 9036 -3385 9052 -3351
rect 10128 -3385 10144 -3351
rect 8790 -3440 8926 -3403
rect 10314 -3403 10341 -2617
rect 10280 -3440 10341 -3403
rect 8790 -3465 10341 -3440
rect 8790 -3499 8962 -3465
rect 10218 -3499 10341 -3465
rect 8790 -3519 10341 -3499
rect 10552 -2507 11179 -2503
rect 12437 -2473 12443 -2335
rect 12477 -2473 12508 -2335
rect 12437 -2507 12508 -2473
rect 10552 -2535 12508 -2507
rect 10552 -2569 11241 -2535
rect 12381 -2569 12508 -2535
rect 10552 -2570 12508 -2569
rect 8679 -3760 10341 -3758
rect 8443 -3769 10341 -3760
rect 10552 -3769 10596 -2570
rect 10669 -2571 12508 -2570
rect 8443 -3820 10596 -3769
rect 3640 -7906 4010 -7895
rect 3586 -7947 4010 -7906
rect 3052 -7968 4010 -7947
rect 3052 -8002 3170 -7968
rect 3544 -8002 4010 -7968
rect 3052 -8023 4010 -8002
rect 3054 -8025 4010 -8023
rect 2313 -8325 2984 -8311
rect 1492 -8337 2984 -8325
rect 1492 -8371 2284 -8337
rect 2866 -8371 2984 -8337
rect 3578 -8356 4010 -8025
rect 3578 -8357 3815 -8356
rect 3578 -8368 3637 -8357
rect 1492 -8418 2984 -8371
rect 3083 -8417 3166 -8368
rect 3545 -8417 3637 -8368
rect 1492 -8423 2105 -8418
rect 1492 -8993 1628 -8423
rect 3083 -8479 3131 -8417
rect 3578 -8444 3637 -8417
rect 3253 -8518 3269 -8484
rect 3445 -8518 3461 -8484
rect 3578 -8486 3602 -8444
rect 3176 -8546 3210 -8530
rect 3176 -8730 3210 -8714
rect 3504 -8546 3538 -8530
rect 3504 -8730 3538 -8714
rect 1492 -9026 2910 -8993
rect 1492 -9060 1680 -9026
rect 1714 -9060 1770 -9026
rect 1804 -9060 1860 -9026
rect 1894 -9060 1950 -9026
rect 1984 -9060 2040 -9026
rect 2074 -9060 2130 -9026
rect 2164 -9060 2220 -9026
rect 2254 -9060 2310 -9026
rect 2344 -9060 2400 -9026
rect 2434 -9060 2490 -9026
rect 2524 -9060 2580 -9026
rect 2614 -9060 2670 -9026
rect 2704 -9060 2760 -9026
rect 2794 -9060 2910 -9026
rect 1492 -9069 2910 -9060
rect 1492 -9127 1720 -9069
rect 1492 -9161 1657 -9127
rect 1691 -9161 1720 -9127
rect 1492 -9177 1720 -9161
rect 2763 -9127 2910 -9069
rect 2763 -9161 2844 -9127
rect 2878 -9161 2910 -9127
rect 2763 -9177 2910 -9161
rect 1492 -9209 1880 -9177
rect 1914 -9209 1970 -9177
rect 2004 -9209 2060 -9177
rect 2094 -9209 2150 -9177
rect 2184 -9209 2240 -9177
rect 2274 -9209 2330 -9177
rect 2364 -9209 2420 -9177
rect 2454 -9209 2510 -9177
rect 2544 -9209 2600 -9177
rect 2634 -9209 2910 -9177
rect 1492 -9217 2910 -9209
rect 1492 -9251 1657 -9217
rect 1691 -9228 2844 -9217
rect 1691 -9233 1857 -9228
rect 1691 -9251 1804 -9233
rect 1492 -9267 1804 -9251
rect 1838 -9267 1857 -9233
rect 1492 -9307 1857 -9267
rect 2675 -9251 2844 -9228
rect 2878 -9251 2910 -9217
rect 2675 -9267 2910 -9251
rect 1492 -9341 1657 -9307
rect 1691 -9323 1857 -9307
rect 1691 -9341 1804 -9323
rect 1492 -9357 1804 -9341
rect 1838 -9357 1857 -9323
rect 1492 -9397 1857 -9357
rect 1492 -9431 1657 -9397
rect 1691 -9413 1857 -9397
rect 1691 -9431 1804 -9413
rect 1492 -9447 1804 -9431
rect 1838 -9447 1857 -9413
rect 1492 -9487 1857 -9447
rect 1492 -9521 1657 -9487
rect 1691 -9503 1857 -9487
rect 1691 -9521 1804 -9503
rect 1492 -9537 1804 -9521
rect 1838 -9537 1857 -9503
rect 1492 -9551 1857 -9537
rect 1492 -10070 1541 -9551
rect 1405 -10078 1541 -10070
rect 1637 -9577 1857 -9551
rect 1637 -9611 1657 -9577
rect 1691 -9593 1857 -9577
rect 1691 -9611 1804 -9593
rect 1637 -9627 1804 -9611
rect 1838 -9627 1857 -9593
rect 1637 -9667 1857 -9627
rect 1637 -9701 1657 -9667
rect 1691 -9683 1857 -9667
rect 1691 -9701 1804 -9683
rect 1637 -9717 1804 -9701
rect 1838 -9717 1857 -9683
rect 1637 -9757 1857 -9717
rect 1637 -9791 1657 -9757
rect 1691 -9773 1857 -9757
rect 1691 -9791 1804 -9773
rect 1637 -9807 1804 -9791
rect 1838 -9807 1857 -9773
rect 1637 -9847 1857 -9807
rect 1637 -9881 1657 -9847
rect 1691 -9863 1857 -9847
rect 1691 -9881 1804 -9863
rect 1637 -9897 1804 -9881
rect 1838 -9897 1857 -9863
rect 1637 -9937 1857 -9897
rect 1637 -9971 1657 -9937
rect 1691 -9953 1857 -9937
rect 1691 -9971 1804 -9953
rect 1637 -9987 1804 -9971
rect 1838 -9987 1857 -9953
rect 1919 -9349 2613 -9290
rect 1919 -9383 1978 -9349
rect 2012 -9377 2068 -9349
rect 2040 -9383 2068 -9377
rect 2102 -9377 2158 -9349
rect 2102 -9383 2106 -9377
rect 1919 -9411 2006 -9383
rect 2040 -9411 2106 -9383
rect 2140 -9383 2158 -9377
rect 2192 -9377 2248 -9349
rect 2192 -9383 2206 -9377
rect 2140 -9411 2206 -9383
rect 2240 -9383 2248 -9377
rect 2282 -9377 2338 -9349
rect 2372 -9377 2428 -9349
rect 2462 -9377 2518 -9349
rect 2282 -9383 2306 -9377
rect 2372 -9383 2406 -9377
rect 2462 -9383 2506 -9377
rect 2552 -9383 2613 -9349
rect 2240 -9411 2306 -9383
rect 2340 -9411 2406 -9383
rect 2440 -9411 2506 -9383
rect 2540 -9411 2613 -9383
rect 1919 -9439 2613 -9411
rect 1919 -9473 1978 -9439
rect 2012 -9473 2068 -9439
rect 2102 -9473 2158 -9439
rect 2192 -9473 2248 -9439
rect 2282 -9473 2338 -9439
rect 2372 -9473 2428 -9439
rect 2462 -9473 2518 -9439
rect 2552 -9473 2613 -9439
rect 1919 -9477 2613 -9473
rect 1919 -9511 2006 -9477
rect 2040 -9511 2106 -9477
rect 2140 -9511 2206 -9477
rect 2240 -9511 2306 -9477
rect 2340 -9511 2406 -9477
rect 2440 -9511 2506 -9477
rect 2540 -9511 2613 -9477
rect 1919 -9529 2613 -9511
rect 1919 -9563 1978 -9529
rect 2012 -9563 2068 -9529
rect 2102 -9563 2158 -9529
rect 2192 -9563 2248 -9529
rect 2282 -9563 2338 -9529
rect 2372 -9563 2428 -9529
rect 2462 -9563 2518 -9529
rect 2552 -9563 2613 -9529
rect 1919 -9577 2613 -9563
rect 1919 -9611 2006 -9577
rect 2040 -9611 2106 -9577
rect 2140 -9611 2206 -9577
rect 2240 -9611 2306 -9577
rect 2340 -9611 2406 -9577
rect 2440 -9611 2506 -9577
rect 2540 -9611 2613 -9577
rect 1919 -9619 2613 -9611
rect 1919 -9653 1978 -9619
rect 2012 -9653 2068 -9619
rect 2102 -9653 2158 -9619
rect 2192 -9653 2248 -9619
rect 2282 -9653 2338 -9619
rect 2372 -9653 2428 -9619
rect 2462 -9653 2518 -9619
rect 2552 -9653 2613 -9619
rect 1919 -9677 2613 -9653
rect 1919 -9709 2006 -9677
rect 2040 -9709 2106 -9677
rect 1919 -9743 1978 -9709
rect 2040 -9711 2068 -9709
rect 2012 -9743 2068 -9711
rect 2102 -9711 2106 -9709
rect 2140 -9709 2206 -9677
rect 2140 -9711 2158 -9709
rect 2102 -9743 2158 -9711
rect 2192 -9711 2206 -9709
rect 2240 -9709 2306 -9677
rect 2340 -9709 2406 -9677
rect 2440 -9709 2506 -9677
rect 2540 -9709 2613 -9677
rect 2240 -9711 2248 -9709
rect 2192 -9743 2248 -9711
rect 2282 -9711 2306 -9709
rect 2372 -9711 2406 -9709
rect 2462 -9711 2506 -9709
rect 2282 -9743 2338 -9711
rect 2372 -9743 2428 -9711
rect 2462 -9743 2518 -9711
rect 2552 -9743 2613 -9709
rect 1919 -9777 2613 -9743
rect 1919 -9799 2006 -9777
rect 2040 -9799 2106 -9777
rect 1919 -9833 1978 -9799
rect 2040 -9811 2068 -9799
rect 2012 -9833 2068 -9811
rect 2102 -9811 2106 -9799
rect 2140 -9799 2206 -9777
rect 2140 -9811 2158 -9799
rect 2102 -9833 2158 -9811
rect 2192 -9811 2206 -9799
rect 2240 -9799 2306 -9777
rect 2340 -9799 2406 -9777
rect 2440 -9799 2506 -9777
rect 2540 -9799 2613 -9777
rect 2240 -9811 2248 -9799
rect 2192 -9833 2248 -9811
rect 2282 -9811 2306 -9799
rect 2372 -9811 2406 -9799
rect 2462 -9811 2506 -9799
rect 2282 -9833 2338 -9811
rect 2372 -9833 2428 -9811
rect 2462 -9833 2518 -9811
rect 2552 -9833 2613 -9799
rect 1919 -9877 2613 -9833
rect 1919 -9889 2006 -9877
rect 2040 -9889 2106 -9877
rect 1919 -9923 1978 -9889
rect 2040 -9911 2068 -9889
rect 2012 -9923 2068 -9911
rect 2102 -9911 2106 -9889
rect 2140 -9889 2206 -9877
rect 2140 -9911 2158 -9889
rect 2102 -9923 2158 -9911
rect 2192 -9911 2206 -9889
rect 2240 -9889 2306 -9877
rect 2340 -9889 2406 -9877
rect 2440 -9889 2506 -9877
rect 2540 -9889 2613 -9877
rect 2240 -9911 2248 -9889
rect 2192 -9923 2248 -9911
rect 2282 -9911 2306 -9889
rect 2372 -9911 2406 -9889
rect 2462 -9911 2506 -9889
rect 2282 -9923 2338 -9911
rect 2372 -9923 2428 -9911
rect 2462 -9923 2518 -9911
rect 2552 -9923 2613 -9889
rect 1919 -9984 2613 -9923
rect 2675 -9301 2694 -9267
rect 2728 -9301 2910 -9267
rect 2675 -9302 2910 -9301
rect 2675 -9357 2730 -9302
rect 2675 -9391 2694 -9357
rect 2728 -9391 2730 -9357
rect 2675 -9447 2730 -9391
rect 2675 -9481 2694 -9447
rect 2728 -9481 2730 -9447
rect 2675 -9537 2730 -9481
rect 2675 -9571 2694 -9537
rect 2728 -9571 2730 -9537
rect 2675 -9627 2730 -9571
rect 2675 -9661 2694 -9627
rect 2728 -9661 2730 -9627
rect 2675 -9717 2730 -9661
rect 2675 -9751 2694 -9717
rect 2728 -9751 2730 -9717
rect 2675 -9807 2730 -9751
rect 2675 -9841 2694 -9807
rect 2728 -9841 2730 -9807
rect 2675 -9897 2730 -9841
rect 2675 -9931 2694 -9897
rect 2728 -9931 2730 -9897
rect 1637 -10027 1857 -9987
rect 1637 -10061 1657 -10027
rect 1691 -10046 1857 -10027
rect 2675 -9987 2730 -9931
rect 2675 -10021 2694 -9987
rect 2728 -10021 2730 -9987
rect 2675 -10046 2730 -10021
rect 1691 -10061 2730 -10046
rect 1637 -10065 2730 -10061
rect 1637 -10078 1861 -10065
rect 1405 -10099 1861 -10078
rect 1895 -10099 1951 -10065
rect 1985 -10099 2041 -10065
rect 2075 -10099 2131 -10065
rect 2165 -10099 2221 -10065
rect 2255 -10099 2311 -10065
rect 2345 -10099 2401 -10065
rect 2435 -10099 2491 -10065
rect 2525 -10099 2581 -10065
rect 2615 -10099 2730 -10065
rect 1405 -10104 2730 -10099
rect 1405 -10117 2153 -10104
rect 1405 -10151 1657 -10117
rect 1691 -10151 2153 -10117
rect 1405 -10187 2153 -10151
rect -1387 -10206 2153 -10187
rect -1387 -10213 -1305 -10206
rect -1153 -10213 -315 -10206
rect -167 -10213 2153 -10206
rect 2632 -10127 2730 -10104
rect 2632 -10151 2844 -10127
rect 2878 -10151 2910 -9302
rect 2632 -10213 2910 -10151
rect -1387 -10247 -1364 -10213
rect 1345 -10247 1680 -10213
rect 1714 -10247 1770 -10213
rect 1804 -10247 1860 -10213
rect 1894 -10247 1950 -10213
rect 1984 -10247 2040 -10213
rect 2074 -10247 2130 -10213
rect 2632 -10224 2670 -10213
rect 2164 -10247 2220 -10224
rect 2254 -10247 2310 -10224
rect 2344 -10247 2400 -10224
rect 2434 -10247 2490 -10224
rect 2524 -10247 2580 -10224
rect 2614 -10247 2670 -10224
rect 2704 -10247 2760 -10213
rect 2794 -10247 2910 -10213
rect -1387 -10260 -1305 -10247
rect -1153 -10260 -315 -10247
rect -167 -10260 2910 -10247
rect -1387 -10263 2910 -10260
rect -1639 -10279 2910 -10263
rect -1639 -10366 -1278 -10279
rect 1536 -10280 2910 -10279
rect 1622 -10281 2910 -10280
rect 3083 -9013 3131 -8756
rect 3253 -8776 3269 -8742
rect 3445 -8776 3461 -8742
rect 3176 -8804 3210 -8788
rect 3176 -8988 3210 -8972
rect 3504 -8804 3538 -8788
rect 3504 -8988 3538 -8972
rect 3253 -9034 3269 -9000
rect 3445 -9034 3461 -9000
rect 3578 -9112 3581 -8486
rect 3253 -9243 3269 -9209
rect 3345 -9243 3361 -9209
rect 3176 -9271 3210 -9255
rect 3176 -9655 3210 -9639
rect 3404 -9271 3438 -9255
rect 3404 -9655 3438 -9639
rect 3253 -9701 3269 -9667
rect 3345 -9701 3361 -9667
rect 3176 -9729 3210 -9713
rect 3176 -10113 3210 -10097
rect 3404 -9729 3438 -9713
rect 3404 -10113 3438 -10097
rect 3575 -10100 3581 -9112
rect 3737 -9343 3815 -8357
rect 3083 -10257 3131 -10121
rect 3253 -10159 3269 -10125
rect 3345 -10159 3361 -10125
rect 3576 -10146 3581 -10100
rect 3575 -10161 3581 -10146
rect 3575 -10257 3604 -10161
rect 3083 -10309 3250 -10257
rect 3486 -10309 3604 -10257
rect 3575 -10336 3604 -10309
rect 3736 -10335 3815 -9343
rect 3963 -8460 4010 -8356
rect 3963 -10335 4009 -8460
rect 3736 -10336 4009 -10335
rect 3575 -10386 4009 -10336
<< viali >>
rect -10213 5416 -2415 5505
rect -9886 5114 -6318 5148
rect -6228 5114 -2660 5148
rect -9948 4719 -9914 5055
rect -6290 4719 -6256 5055
rect -2632 4719 -2598 5055
rect -9886 4626 -6318 4660
rect -6228 4626 -2660 4660
rect -9948 4231 -9914 4567
rect -6290 4231 -6256 4567
rect -2632 4231 -2598 4567
rect -9886 4138 -6318 4172
rect -6228 4138 -2660 4172
rect -1814 7557 778 7627
rect -1814 7523 -1680 7557
rect -1680 7523 600 7557
rect 600 7523 778 7557
rect -1814 7497 778 7523
rect -1814 4016 -1740 7497
rect -1740 4016 -1706 7497
rect -1706 7424 626 7497
rect 626 7424 660 7497
rect 660 7424 778 7497
rect -1706 4016 -1649 7424
rect -1414 7190 -1066 7224
rect -976 7190 -628 7224
rect -538 7190 -190 7224
rect -100 7190 248 7224
rect -1476 4155 -1442 7131
rect -1038 4155 -1004 7131
rect -600 4155 -566 7131
rect -162 4155 -128 7131
rect 276 4155 310 7131
rect 566 4365 626 6845
rect 626 4365 660 6845
rect 660 4365 708 6845
rect -1414 4062 -1066 4096
rect -976 4062 -628 4096
rect -538 4062 -190 4096
rect -100 4062 248 4096
rect -10065 1636 -9489 1670
rect -10149 640 -10115 1608
rect -9439 640 -9405 1608
rect -10065 578 -9489 612
rect -10291 -26 -9738 68
rect -8676 3233 -6308 3267
rect -6218 3233 -3850 3267
rect -8738 2007 -8704 3183
rect -6280 2007 -6246 3183
rect -3822 2007 -3788 3183
rect -8676 1923 -6308 1957
rect -6218 1923 -3850 1957
rect -8677 1358 -6309 1392
rect -6219 1358 -3851 1392
rect -8739 132 -8705 1308
rect -6281 132 -6247 1308
rect -3823 132 -3789 1308
rect -8677 48 -6309 82
rect -6219 48 -3851 82
rect -1414 3213 -1066 3247
rect -976 3213 -628 3247
rect -538 3213 -190 3247
rect -100 3213 248 3247
rect -1797 22 -1740 3198
rect -1798 -38 -1740 22
rect -1740 -38 -1706 3198
rect -1706 -11 -1649 3198
rect -1476 178 -1442 3154
rect -1038 178 -1004 3154
rect -600 178 -566 3154
rect -162 178 -128 3154
rect 276 178 310 3154
rect 582 132 626 2612
rect 626 132 660 2612
rect 660 2114 724 2612
rect 11789 2772 12048 2773
rect 7086 2473 12048 2772
rect 7086 2439 7241 2473
rect 7241 2439 11927 2473
rect 11927 2439 12048 2473
rect 7086 2413 12048 2439
rect 7086 2407 7181 2413
rect 660 2113 5514 2114
rect 660 1822 5524 2113
rect 660 132 724 1822
rect -1414 85 -1066 119
rect -976 85 -628 119
rect -538 85 -190 119
rect -100 85 248 119
rect -1706 -38 626 -11
rect 626 -38 660 -11
rect 660 -38 767 -11
rect -1798 -64 767 -38
rect -1798 -98 -1680 -64
rect -1680 -98 600 -64
rect 600 -98 767 -64
rect -1798 -154 767 -98
rect -1685 -155 767 -154
rect -10289 -256 -3355 -167
rect 2986 66 3219 1822
rect 3415 1659 3743 1693
rect 3833 1659 4161 1693
rect 4251 1659 4579 1693
rect 4669 1659 4997 1693
rect 3353 224 3387 1600
rect 3771 224 3805 1600
rect 4189 224 4223 1600
rect 4607 224 4641 1600
rect 5025 224 5059 1600
rect 3415 131 3743 165
rect 3833 131 4161 165
rect 4251 131 4579 165
rect 4669 131 4997 165
rect 5237 306 5524 1822
rect 7148 200 7181 2407
rect 7181 200 7215 2413
rect 7215 2408 11953 2413
rect 7215 2407 11890 2408
rect 7215 205 7265 2407
rect 7508 2204 8476 2238
rect 8566 2204 9534 2238
rect 9624 2204 10592 2238
rect 10682 2204 11650 2238
rect 7446 1669 7480 2145
rect 8504 1669 8538 2145
rect 9562 1669 9596 2145
rect 10620 1669 10654 2145
rect 11678 1669 11712 2145
rect 7508 1576 8476 1610
rect 8566 1576 9534 1610
rect 9624 1576 10592 1610
rect 10682 1576 11650 1610
rect 11932 1594 11953 2408
rect 11953 1594 11987 2413
rect 11987 2408 12048 2413
rect 11987 1594 12029 2408
rect 7508 1042 8476 1076
rect 8566 1042 9534 1076
rect 9624 1042 10592 1076
rect 10682 1042 11650 1076
rect 7446 507 7480 983
rect 8504 507 8538 983
rect 9562 507 9596 983
rect 10620 507 10654 983
rect 11678 507 11712 983
rect 7508 414 8476 448
rect 8566 414 9534 448
rect 9624 414 10592 448
rect 10682 414 11650 448
rect 7215 200 11697 205
rect 7148 174 11697 200
rect 7148 140 7241 174
rect 7241 140 11697 174
rect 7148 115 11697 140
rect 7183 108 11697 115
rect 2986 63 5134 66
rect 2986 29 3335 63
rect 3335 29 5077 63
rect 5077 29 5134 63
rect 2986 -168 5134 29
rect 3071 -170 5134 -168
rect 8506 -74 10655 -25
rect 8506 -108 8581 -74
rect 8581 -108 10563 -74
rect 10563 -108 10655 -74
rect 8506 -128 10655 -108
rect 8506 -134 8564 -128
rect -1742 -496 -1595 -493
rect 6084 -496 6200 -456
rect -1742 -530 -1628 -496
rect -1628 -501 -1595 -496
rect -1628 -502 -1466 -501
rect 6084 -502 6200 -496
rect -1628 -530 6200 -502
rect -1742 -556 6200 -530
rect -1742 -1779 -1688 -556
rect -1688 -1779 -1654 -556
rect -1654 -605 6200 -556
rect -1654 -1779 -1595 -605
rect 6084 -617 6200 -605
rect -1404 -822 444 -788
rect 534 -822 2382 -788
rect 2472 -822 4320 -788
rect 4410 -822 6258 -788
rect -1466 -1148 -1432 -872
rect 472 -1148 506 -872
rect 2410 -1148 2444 -872
rect 4348 -1148 4382 -872
rect 6286 -1148 6320 -872
rect -1404 -1232 444 -1198
rect 534 -1232 2382 -1198
rect 2472 -1232 4320 -1198
rect 4410 -1232 6258 -1198
rect -1466 -1558 -1432 -1282
rect 472 -1558 506 -1282
rect 2410 -1558 2444 -1282
rect 4348 -1558 4382 -1282
rect 6286 -1558 6320 -1282
rect -1404 -1642 444 -1608
rect 534 -1642 2382 -1608
rect 2472 -1642 4320 -1608
rect 4410 -1642 6258 -1608
rect -1742 -1795 -1595 -1779
rect -1742 -1796 -1501 -1795
rect -1742 -1805 6177 -1796
rect -1742 -1839 -1628 -1805
rect -1628 -1839 6177 -1805
rect -1742 -1993 6177 -1839
rect 8506 -666 8521 -134
rect 8521 -666 8555 -134
rect 8555 -666 8564 -134
rect 10579 -134 10655 -128
rect 8693 -252 9061 -218
rect 9151 -252 9519 -218
rect 9609 -252 9977 -218
rect 10067 -252 10435 -218
rect 8631 -878 8665 -302
rect 9089 -878 9123 -302
rect 9547 -878 9581 -302
rect 10005 -878 10039 -302
rect 10463 -878 10497 -302
rect 8693 -962 9061 -928
rect 9151 -962 9519 -928
rect 9609 -962 9977 -928
rect 10067 -962 10435 -928
rect 8693 -1459 9061 -1425
rect 9151 -1459 9519 -1425
rect 9609 -1459 9977 -1425
rect 10067 -1459 10435 -1425
rect 8497 -2252 8521 -1702
rect 8521 -2252 8555 -1702
rect 8555 -2252 8571 -1702
rect 8631 -2085 8665 -1509
rect 9089 -2085 9123 -1509
rect 9547 -2085 9581 -1509
rect 10005 -2085 10039 -1509
rect 10463 -2085 10497 -1509
rect 8693 -2169 9061 -2135
rect 9151 -2169 9519 -2135
rect 9609 -2169 9977 -2135
rect 10067 -2169 10435 -2135
rect 8497 -2333 8571 -2252
rect 10579 -2252 10589 -134
rect 10589 -2252 10623 -134
rect 10623 -2252 10655 -134
rect 11593 -321 11697 108
rect 11593 -1015 11665 -321
rect 11665 -1015 11697 -321
rect 11841 -361 11879 -327
rect 11779 -916 11813 -420
rect 11907 -916 11941 -420
rect 11841 -1009 11879 -975
rect 11593 -1051 11697 -1015
rect 12197 -361 12235 -327
rect 12135 -916 12169 -420
rect 12263 -916 12297 -420
rect 12197 -1009 12235 -975
rect 11863 -1375 11897 -1341
rect 12219 -1375 12253 -1341
rect 11819 -1601 11853 -1425
rect 11907 -1601 11941 -1425
rect 12175 -1601 12209 -1425
rect 12263 -1601 12297 -1425
rect 11863 -1685 11897 -1651
rect 12219 -1685 12253 -1651
rect 10997 -2157 12375 -1885
rect 10579 -2333 10655 -2252
rect 10997 -2333 11117 -2157
rect 8452 -2503 11117 -2333
rect 11293 -2423 11690 -2385
rect 11932 -2423 12329 -2385
rect -1561 -3731 -1387 -3685
rect 1380 -3731 1492 -3729
rect -1561 -10187 -1424 -3731
rect -1424 -10187 -1390 -3731
rect -1390 -10187 -1387 -3731
rect -1136 -3849 -360 -3815
rect 345 -3849 1121 -3815
rect -1220 -4045 -1186 -3877
rect -310 -4045 -276 -3877
rect 261 -4045 295 -3877
rect 1171 -4045 1205 -3877
rect -1136 -4107 -360 -4073
rect 345 -4107 1121 -4073
rect -1220 -4303 -1186 -4135
rect -310 -4303 -276 -4135
rect 261 -4303 295 -4135
rect 1171 -4303 1205 -4135
rect -1136 -4365 -360 -4331
rect 345 -4365 1121 -4331
rect -1220 -4561 -1186 -4393
rect -310 -4561 -276 -4393
rect 261 -4561 295 -4393
rect 1171 -4561 1205 -4393
rect -1136 -4623 -360 -4589
rect 345 -4623 1121 -4589
rect -1220 -4819 -1186 -4651
rect -310 -4819 -276 -4651
rect 261 -4819 295 -4651
rect 1171 -4819 1205 -4651
rect -1136 -4881 -360 -4847
rect 345 -4881 1121 -4847
rect -1220 -5077 -1186 -4909
rect -310 -5077 -276 -4909
rect 261 -5077 295 -4909
rect 1171 -5077 1205 -4909
rect -1136 -5139 -360 -5105
rect 345 -5139 1121 -5105
rect -1220 -5335 -1186 -5167
rect -310 -5335 -276 -5167
rect 261 -5335 295 -5167
rect 1171 -5335 1205 -5167
rect -1136 -5397 -360 -5363
rect 345 -5397 1121 -5363
rect -1220 -5593 -1186 -5425
rect -310 -5593 -276 -5425
rect 261 -5593 295 -5425
rect 1171 -5593 1205 -5425
rect -1136 -5655 -360 -5621
rect 345 -5655 1121 -5621
rect -1220 -5851 -1186 -5683
rect -310 -5851 -276 -5683
rect 261 -5851 295 -5683
rect 1171 -5851 1205 -5683
rect -1136 -5913 -360 -5879
rect 345 -5913 1121 -5879
rect -1220 -6109 -1186 -5941
rect -310 -6109 -276 -5941
rect 261 -6109 295 -5941
rect 1171 -6109 1205 -5941
rect -1136 -6171 -360 -6137
rect 345 -6171 1121 -6137
rect -1220 -6367 -1186 -6199
rect -310 -6367 -276 -6199
rect 261 -6367 295 -6199
rect 1171 -6367 1205 -6199
rect -1136 -6429 -360 -6395
rect 345 -6429 1121 -6395
rect -1220 -6625 -1186 -6457
rect -310 -6625 -276 -6457
rect 261 -6625 295 -6457
rect 1171 -6625 1205 -6457
rect -1136 -6687 -360 -6653
rect 345 -6687 1121 -6653
rect -1220 -6883 -1186 -6715
rect -310 -6883 -276 -6715
rect 261 -6883 295 -6715
rect 1171 -6883 1205 -6715
rect -1136 -6945 -360 -6911
rect 345 -6945 1121 -6911
rect -1220 -7141 -1186 -6973
rect -310 -7141 -276 -6973
rect 261 -7141 295 -6973
rect 1171 -7141 1205 -6973
rect -1136 -7203 -360 -7169
rect 345 -7203 1121 -7169
rect -1220 -7399 -1186 -7231
rect -310 -7399 -276 -7231
rect 261 -7399 295 -7231
rect 1171 -7399 1205 -7231
rect -1136 -7461 -360 -7427
rect 345 -7461 1121 -7427
rect -1220 -7657 -1186 -7489
rect -310 -7657 -276 -7489
rect 261 -7657 295 -7489
rect 1171 -7657 1205 -7489
rect -1136 -7719 -360 -7685
rect 345 -7719 1121 -7685
rect -1220 -7915 -1186 -7747
rect -310 -7915 -276 -7747
rect 261 -7915 295 -7747
rect 1171 -7915 1205 -7747
rect -1136 -7977 -360 -7943
rect 345 -7977 1121 -7943
rect -1220 -8173 -1186 -8005
rect -310 -8173 -276 -8005
rect 261 -8173 295 -8005
rect 1171 -8173 1205 -8005
rect -1136 -8235 -360 -8201
rect 345 -8235 1121 -8201
rect -1220 -8431 -1186 -8263
rect -310 -8431 -276 -8263
rect 261 -8431 295 -8263
rect 1171 -8431 1205 -8263
rect -1136 -8493 -360 -8459
rect 345 -8493 1121 -8459
rect -1220 -8689 -1186 -8521
rect -310 -8689 -276 -8521
rect 261 -8689 295 -8521
rect 1171 -8689 1205 -8521
rect -1136 -8751 -360 -8717
rect 345 -8751 1121 -8717
rect -1220 -8947 -1186 -8779
rect -310 -8947 -276 -8779
rect 261 -8947 295 -8779
rect 1171 -8947 1205 -8779
rect -1136 -9009 -360 -8975
rect 345 -9009 1121 -8975
rect -1220 -9205 -1186 -9037
rect -310 -9205 -276 -9037
rect 261 -9205 295 -9037
rect 1171 -9205 1205 -9037
rect -1136 -9267 -360 -9233
rect 345 -9267 1121 -9233
rect -1220 -9463 -1186 -9295
rect -310 -9463 -276 -9295
rect 261 -9463 295 -9295
rect 1171 -9463 1205 -9295
rect -1136 -9525 -360 -9491
rect 345 -9525 1121 -9491
rect -1220 -9721 -1186 -9553
rect -310 -9721 -276 -9553
rect 261 -9721 295 -9553
rect 1171 -9721 1205 -9553
rect -1136 -9783 -360 -9749
rect 345 -9783 1121 -9749
rect -1220 -9979 -1186 -9811
rect -310 -9979 -276 -9811
rect 261 -9979 295 -9811
rect 1171 -9979 1205 -9811
rect -1136 -10041 -360 -10007
rect 345 -10041 1121 -10007
rect 1380 -10070 1405 -3731
rect 1405 -10070 1492 -3731
rect 2122 -8311 2224 -2918
rect 2224 -8311 2258 -2918
rect 2258 -8311 2313 -2918
rect 2482 -3044 2658 -3010
rect 2398 -3240 2432 -3072
rect 2708 -3240 2742 -3072
rect 2482 -3302 2658 -3268
rect 2398 -3498 2432 -3330
rect 2708 -3498 2742 -3330
rect 2482 -3560 2658 -3526
rect 2398 -3756 2432 -3588
rect 2708 -3756 2742 -3588
rect 2482 -3818 2658 -3784
rect 2398 -4014 2432 -3846
rect 2708 -4014 2742 -3846
rect 2482 -4076 2658 -4042
rect 2398 -4272 2432 -4104
rect 2708 -4272 2742 -4104
rect 2482 -4334 2658 -4300
rect 2398 -4530 2432 -4362
rect 2708 -4530 2742 -4362
rect 2482 -4592 2658 -4558
rect 2398 -4788 2432 -4620
rect 2708 -4788 2742 -4620
rect 2482 -4850 2658 -4816
rect 2398 -5046 2432 -4878
rect 2708 -5046 2742 -4878
rect 2482 -5108 2658 -5074
rect 2398 -5304 2432 -5136
rect 2708 -5304 2742 -5136
rect 2482 -5366 2658 -5332
rect 2398 -5562 2432 -5394
rect 2708 -5562 2742 -5394
rect 2482 -5624 2658 -5590
rect 2398 -5820 2432 -5652
rect 2708 -5820 2742 -5652
rect 2482 -5882 2658 -5848
rect 2398 -6078 2432 -5910
rect 2708 -6078 2742 -5910
rect 2482 -6140 2658 -6106
rect 2398 -6336 2432 -6168
rect 2708 -6336 2742 -6168
rect 2482 -6398 2658 -6364
rect 2398 -6594 2432 -6426
rect 2708 -6594 2742 -6426
rect 2482 -6656 2658 -6622
rect 2398 -6852 2432 -6684
rect 2708 -6852 2742 -6684
rect 2482 -6914 2658 -6880
rect 2398 -7110 2432 -6942
rect 2708 -7110 2742 -6942
rect 2482 -7172 2658 -7138
rect 2398 -7368 2432 -7200
rect 2708 -7368 2742 -7200
rect 2482 -7430 2658 -7396
rect 2398 -7626 2432 -7458
rect 2708 -7626 2742 -7458
rect 2482 -7688 2658 -7654
rect 2398 -7884 2432 -7716
rect 2708 -7884 2742 -7716
rect 2482 -7946 2658 -7912
rect 2398 -8142 2432 -7974
rect 2708 -8142 2742 -7974
rect 2482 -8204 2658 -8170
rect 3269 -2979 3445 -2945
rect 3176 -3375 3210 -3007
rect 3504 -3375 3538 -3007
rect 3269 -3437 3445 -3403
rect 3269 -3560 3445 -3526
rect 3176 -3956 3210 -3588
rect 3504 -3956 3538 -3588
rect 3269 -4018 3445 -3984
rect 3269 -4850 3445 -4816
rect 3176 -5246 3210 -4878
rect 3504 -5246 3538 -4878
rect 3269 -5308 3445 -5274
rect 3269 -6140 3445 -6106
rect 3176 -6536 3210 -6168
rect 3504 -6536 3538 -6168
rect 3269 -6598 3445 -6564
rect 3269 -7430 3445 -7396
rect 3176 -7826 3210 -7458
rect 3504 -7826 3538 -7458
rect 3269 -7888 3445 -7854
rect 3716 -7895 3855 -2900
rect 8452 -3519 8790 -2503
rect 9052 -2669 10128 -2635
rect 8968 -2965 9002 -2697
rect 10178 -2965 10212 -2697
rect 9052 -3027 10128 -2993
rect 8968 -3323 9002 -3055
rect 10178 -3323 10212 -3055
rect 9052 -3385 10128 -3351
rect 10341 -3519 10552 -2503
rect 8452 -3758 10552 -3519
rect 8452 -3760 8679 -3758
rect 10341 -3769 10552 -3758
rect 2122 -8325 2313 -8311
rect 3637 -8444 3737 -8357
rect 3269 -8518 3445 -8484
rect 3602 -8486 3737 -8444
rect 3176 -8714 3210 -8546
rect 3504 -8714 3538 -8546
rect 1720 -9175 2763 -9069
rect 1720 -9177 1880 -9175
rect 1880 -9177 1914 -9175
rect 1914 -9177 1970 -9175
rect 1970 -9177 2004 -9175
rect 2004 -9177 2060 -9175
rect 2060 -9177 2094 -9175
rect 2094 -9177 2150 -9175
rect 2150 -9177 2184 -9175
rect 2184 -9177 2240 -9175
rect 2240 -9177 2274 -9175
rect 2274 -9177 2330 -9175
rect 2330 -9177 2364 -9175
rect 2364 -9177 2420 -9175
rect 2420 -9177 2454 -9175
rect 2454 -9177 2510 -9175
rect 2510 -9177 2544 -9175
rect 2544 -9177 2600 -9175
rect 2600 -9177 2634 -9175
rect 2634 -9177 2763 -9175
rect 1541 -10078 1637 -9551
rect 2006 -9383 2012 -9377
rect 2012 -9383 2040 -9377
rect 2006 -9411 2040 -9383
rect 2106 -9411 2140 -9377
rect 2206 -9411 2240 -9377
rect 2306 -9383 2338 -9377
rect 2338 -9383 2340 -9377
rect 2406 -9383 2428 -9377
rect 2428 -9383 2440 -9377
rect 2506 -9383 2518 -9377
rect 2518 -9383 2540 -9377
rect 2306 -9411 2340 -9383
rect 2406 -9411 2440 -9383
rect 2506 -9411 2540 -9383
rect 2006 -9511 2040 -9477
rect 2106 -9511 2140 -9477
rect 2206 -9511 2240 -9477
rect 2306 -9511 2340 -9477
rect 2406 -9511 2440 -9477
rect 2506 -9511 2540 -9477
rect 2006 -9611 2040 -9577
rect 2106 -9611 2140 -9577
rect 2206 -9611 2240 -9577
rect 2306 -9611 2340 -9577
rect 2406 -9611 2440 -9577
rect 2506 -9611 2540 -9577
rect 2006 -9709 2040 -9677
rect 2006 -9711 2012 -9709
rect 2012 -9711 2040 -9709
rect 2106 -9711 2140 -9677
rect 2206 -9711 2240 -9677
rect 2306 -9709 2340 -9677
rect 2406 -9709 2440 -9677
rect 2506 -9709 2540 -9677
rect 2306 -9711 2338 -9709
rect 2338 -9711 2340 -9709
rect 2406 -9711 2428 -9709
rect 2428 -9711 2440 -9709
rect 2506 -9711 2518 -9709
rect 2518 -9711 2540 -9709
rect 2006 -9799 2040 -9777
rect 2006 -9811 2012 -9799
rect 2012 -9811 2040 -9799
rect 2106 -9811 2140 -9777
rect 2206 -9811 2240 -9777
rect 2306 -9799 2340 -9777
rect 2406 -9799 2440 -9777
rect 2506 -9799 2540 -9777
rect 2306 -9811 2338 -9799
rect 2338 -9811 2340 -9799
rect 2406 -9811 2428 -9799
rect 2428 -9811 2440 -9799
rect 2506 -9811 2518 -9799
rect 2518 -9811 2540 -9799
rect 2006 -9889 2040 -9877
rect 2006 -9911 2012 -9889
rect 2012 -9911 2040 -9889
rect 2106 -9911 2140 -9877
rect 2206 -9911 2240 -9877
rect 2306 -9889 2340 -9877
rect 2406 -9889 2440 -9877
rect 2506 -9889 2540 -9877
rect 2306 -9911 2338 -9889
rect 2338 -9911 2340 -9889
rect 2406 -9911 2428 -9889
rect 2428 -9911 2440 -9889
rect 2506 -9911 2518 -9889
rect 2518 -9911 2540 -9889
rect 2730 -9307 2878 -9302
rect 2730 -9341 2844 -9307
rect 2844 -9341 2878 -9307
rect 2730 -9397 2878 -9341
rect 2730 -9431 2844 -9397
rect 2844 -9431 2878 -9397
rect 2730 -9487 2878 -9431
rect 2730 -9521 2844 -9487
rect 2844 -9521 2878 -9487
rect 2730 -9577 2878 -9521
rect 2730 -9611 2844 -9577
rect 2844 -9611 2878 -9577
rect 2730 -9667 2878 -9611
rect 2730 -9701 2844 -9667
rect 2844 -9701 2878 -9667
rect 2730 -9757 2878 -9701
rect 2730 -9791 2844 -9757
rect 2844 -9791 2878 -9757
rect 2730 -9847 2878 -9791
rect 2730 -9881 2844 -9847
rect 2844 -9881 2878 -9847
rect 2730 -9937 2878 -9881
rect 2730 -9971 2844 -9937
rect 2844 -9971 2878 -9937
rect 2730 -10027 2878 -9971
rect 2730 -10061 2844 -10027
rect 2844 -10061 2878 -10027
rect -1561 -10263 -1387 -10187
rect -1305 -10213 -1153 -10206
rect -315 -10213 -167 -10206
rect 2153 -10213 2632 -10104
rect 2730 -10117 2878 -10061
rect 2730 -10127 2844 -10117
rect 2844 -10127 2878 -10117
rect -1305 -10247 -1153 -10213
rect -315 -10247 -167 -10213
rect 2153 -10224 2164 -10213
rect 2164 -10224 2220 -10213
rect 2220 -10224 2254 -10213
rect 2254 -10224 2310 -10213
rect 2310 -10224 2344 -10213
rect 2344 -10224 2400 -10213
rect 2400 -10224 2434 -10213
rect 2434 -10224 2490 -10213
rect 2490 -10224 2524 -10213
rect 2524 -10224 2580 -10213
rect 2580 -10224 2614 -10213
rect 2614 -10224 2632 -10213
rect -1305 -10260 -1153 -10247
rect -315 -10260 -167 -10247
rect 3269 -8776 3445 -8742
rect 3176 -8972 3210 -8804
rect 3504 -8972 3538 -8804
rect 3269 -9034 3445 -9000
rect 3269 -9243 3345 -9209
rect 3176 -9639 3210 -9271
rect 3404 -9639 3438 -9271
rect 3269 -9701 3345 -9667
rect 3176 -10097 3210 -9729
rect 3404 -10097 3438 -9729
rect 3602 -9343 3633 -8486
rect 3633 -9343 3737 -8486
rect 3269 -10159 3345 -10125
rect 3604 -10161 3633 -9343
rect 3633 -10161 3736 -9343
rect 3604 -10336 3736 -10161
rect 3815 -10335 3963 -8356
<< metal1 >>
rect -1826 7627 790 7633
rect -1826 7418 -1814 7627
rect 778 7424 790 7627
rect -10225 5505 -2403 5511
rect -10225 5416 -10213 5505
rect -2415 5416 -2403 5505
rect -10225 5410 -2403 5416
rect -10095 5148 -2648 5154
rect -10095 5114 -9886 5148
rect -6318 5114 -6228 5148
rect -2660 5114 -2648 5148
rect -10095 5108 -2648 5114
rect -10095 5055 -9895 5108
rect -10095 4719 -9948 5055
rect -9914 4719 -9895 5055
rect -10095 4706 -9895 4719
rect -10095 3675 -10009 4706
rect -9718 4666 -6479 5108
rect -6296 5055 -6250 5067
rect -6310 4719 -6300 5055
rect -6246 4719 -6236 5055
rect -6296 4707 -6250 4719
rect -6056 4666 -2817 5108
rect -2652 5055 -2450 5068
rect -2652 4719 -2632 5055
rect -2598 4719 -2450 5055
rect -2652 4708 -2450 4719
rect -2638 4707 -2592 4708
rect -9898 4660 -6306 4666
rect -9898 4626 -9886 4660
rect -6318 4626 -6306 4660
rect -9898 4620 -6306 4626
rect -6240 4660 -2648 4666
rect -6240 4626 -6228 4660
rect -2660 4626 -2648 4660
rect -6240 4620 -2648 4626
rect -9981 4567 -9895 4579
rect -9981 4536 -9948 4567
rect -9914 4536 -9895 4567
rect -9905 4231 -9895 4536
rect -9981 4218 -9895 4231
rect -9718 4178 -6479 4620
rect -6296 4567 -6250 4579
rect -6310 4231 -6300 4567
rect -6246 4231 -6236 4567
rect -6296 4219 -6250 4231
rect -6056 4178 -2817 4620
rect -2650 4567 -2564 4579
rect -2650 4526 -2632 4567
rect -2598 4526 -2564 4567
rect -2650 4231 -2640 4526
rect -2650 4178 -2564 4231
rect -9898 4172 -2564 4178
rect -9898 4138 -9886 4172
rect -6318 4138 -6228 4172
rect -2660 4138 -2564 4172
rect -9898 4132 -2564 4138
rect -2536 3860 -2450 4708
rect -1824 4016 -1814 7418
rect -1649 7418 790 7424
rect -1649 4016 -1639 7418
rect -1426 7224 -1054 7230
rect -1426 7190 -1414 7224
rect -1066 7190 -1054 7224
rect -1426 7184 -1054 7190
rect -988 7224 -616 7230
rect -988 7190 -976 7224
rect -628 7190 -616 7224
rect -988 7184 -616 7190
rect -550 7224 -178 7230
rect -550 7190 -538 7224
rect -190 7190 -178 7224
rect -550 7184 -178 7190
rect -112 7224 260 7230
rect -112 7190 -100 7224
rect 248 7190 260 7224
rect -112 7184 260 7190
rect -1482 7131 -1436 7143
rect -1482 5155 -1476 7131
rect -1442 5155 -1436 7131
rect -1502 4155 -1492 5155
rect -1428 4155 -1418 5155
rect -1482 4143 -1436 4155
rect -1354 4105 -1149 7184
rect -1044 7131 -998 7143
rect -1067 6531 -1057 7131
rect -985 6531 -975 7131
rect -1044 4155 -1038 6531
rect -1004 4155 -998 6531
rect -1044 4143 -998 4155
rect -901 4105 -696 7184
rect -606 7131 -560 7143
rect -606 6392 -600 7131
rect -566 6392 -560 7131
rect -625 5392 -615 6392
rect -551 5392 -541 6392
rect -606 4155 -600 5392
rect -566 4155 -560 5392
rect -606 4143 -560 4155
rect -465 4105 -260 7184
rect -168 7131 -122 7143
rect -191 6531 -181 7131
rect -109 6531 -99 7131
rect -168 4155 -162 6531
rect -128 4155 -122 6531
rect -168 4143 -122 4155
rect -25 4105 180 7184
rect 270 7131 316 7143
rect 270 5155 276 7131
rect 310 5155 316 7131
rect 560 6845 714 6857
rect 251 4155 261 5155
rect 325 4155 335 5155
rect 560 4365 566 6845
rect 708 4365 714 6845
rect 560 4353 714 4365
rect 270 4143 316 4155
rect -1424 4102 -1414 4105
rect -1426 4056 -1414 4102
rect -1134 4102 -1124 4105
rect -986 4102 -976 4105
rect -1134 4096 -1054 4102
rect -1066 4062 -1054 4096
rect -1424 4053 -1414 4056
rect -1134 4056 -1054 4062
rect -988 4056 -976 4102
rect -696 4102 -686 4105
rect -548 4102 -538 4105
rect -696 4096 -616 4102
rect -628 4062 -616 4096
rect -1134 4053 -1124 4056
rect -986 4053 -976 4056
rect -696 4056 -616 4062
rect -550 4056 -538 4102
rect -258 4102 -248 4105
rect -110 4102 -100 4105
rect -258 4096 -178 4102
rect -190 4062 -178 4096
rect -696 4053 -686 4056
rect -548 4053 -538 4056
rect -258 4056 -178 4062
rect -112 4056 -100 4102
rect 180 4102 190 4105
rect 180 4096 260 4102
rect 248 4062 260 4096
rect -258 4053 -248 4056
rect -110 4053 -100 4056
rect 180 4056 260 4062
rect 180 4053 190 4056
rect -1820 4004 -1643 4016
rect -9981 3853 -1414 3860
rect -9672 3845 -1414 3853
rect -9672 3778 -9173 3845
rect -8824 3842 -1414 3845
rect -8824 3778 -4109 3842
rect -9672 3775 -4109 3778
rect -3760 3775 -1414 3842
rect -9672 3769 -1414 3775
rect -9981 3760 -1414 3769
rect -1314 3760 -728 3860
rect -628 3760 -290 3860
rect -190 3760 -100 3860
rect 0 3760 1725 3860
rect 2007 3760 2017 3860
rect -10095 3659 -2554 3675
rect -10095 3655 -3689 3659
rect -10095 3588 -8746 3655
rect -8397 3592 -3689 3655
rect -3340 3592 -2975 3659
rect -8397 3589 -2975 3592
rect -2585 3589 -2554 3659
rect -8397 3588 -2554 3589
rect -10095 3575 -2554 3588
rect -2640 3551 -2554 3575
rect -2640 3451 -1166 3551
rect -1066 3451 -976 3551
rect -876 3451 -538 3551
rect -438 3451 148 3551
rect 248 3451 405 3551
rect -8688 3267 -6296 3273
rect -8688 3233 -8676 3267
rect -6308 3233 -6296 3267
rect -8688 3227 -6296 3233
rect -6230 3267 -3838 3273
rect -6230 3233 -6218 3267
rect -3850 3233 -3838 3267
rect -1356 3253 -1346 3256
rect -6230 3227 -3838 3233
rect -1426 3247 -1346 3253
rect -1066 3253 -1056 3256
rect -918 3253 -908 3256
rect -8744 3183 -8698 3195
rect -8792 2615 -8782 3183
rect -8696 2615 -8686 3183
rect -8792 2049 -8738 2615
rect -8744 2007 -8738 2049
rect -8704 2049 -8686 2615
rect -8704 2007 -8698 2049
rect -8744 1995 -8698 2007
rect -8040 1969 -6955 3227
rect -6286 3183 -6240 3195
rect -6286 2358 -6280 3183
rect -6246 2358 -6240 3183
rect -6298 2039 -6288 2358
rect -6236 2039 -6226 2358
rect -6286 2007 -6280 2039
rect -6246 2007 -6240 2039
rect -6286 1995 -6240 2007
rect -5536 1969 -4449 3227
rect -1426 3213 -1414 3247
rect -1803 3198 -1643 3210
rect -1426 3207 -1346 3213
rect -1356 3204 -1346 3207
rect -1066 3207 -1054 3253
rect -988 3247 -908 3253
rect -628 3253 -618 3256
rect -480 3253 -470 3256
rect -988 3213 -976 3247
rect -988 3207 -908 3213
rect -1066 3204 -1056 3207
rect -918 3204 -908 3207
rect -628 3207 -616 3253
rect -550 3247 -470 3253
rect -190 3253 -180 3256
rect -42 3253 -32 3256
rect -550 3213 -538 3247
rect -550 3207 -470 3213
rect -628 3204 -618 3207
rect -480 3204 -470 3207
rect -190 3207 -178 3253
rect -112 3247 -32 3253
rect 248 3253 258 3256
rect -112 3213 -100 3247
rect -112 3207 -32 3213
rect -190 3204 -180 3207
rect -42 3204 -32 3207
rect 248 3207 260 3253
rect 248 3204 258 3207
rect -3828 3183 -3782 3195
rect -3840 2615 -3830 3183
rect -3744 2615 -3734 3183
rect -3840 2062 -3822 2615
rect -3828 2007 -3822 2062
rect -3788 2062 -3734 2615
rect -3788 2007 -3782 2062
rect -3828 1995 -3782 2007
rect -8682 1963 -8672 1969
rect -8688 1957 -8672 1963
rect -8462 1963 -6298 1969
rect -6228 1963 -4060 1969
rect -8462 1957 -6296 1963
rect -8688 1923 -8676 1957
rect -6308 1923 -6296 1957
rect -8688 1917 -8672 1923
rect -8682 1912 -8672 1917
rect -8462 1917 -6296 1923
rect -6230 1957 -4060 1963
rect -3850 1963 -3840 1969
rect -6230 1923 -6218 1957
rect -6230 1917 -4060 1923
rect -8462 1912 -6298 1917
rect -6228 1912 -4060 1917
rect -3850 1917 -3838 1963
rect -3850 1912 -3840 1917
rect -8672 1851 -6219 1855
rect -8672 1794 -8649 1851
rect -8462 1794 -6219 1851
rect -8672 1791 -6219 1794
rect -6018 1791 -6009 1855
rect -8672 1776 -6009 1791
rect -10075 1676 -10065 1687
rect -10077 1632 -10065 1676
rect -9489 1676 -9479 1687
rect -9489 1632 -9477 1676
rect -10077 1630 -9477 1632
rect -10155 1608 -10109 1620
rect -10155 640 -10149 1608
rect -10115 1421 -10109 1608
rect -9445 1608 -9386 1620
rect -9445 1439 -9439 1608
rect -9405 1439 -9386 1608
rect -6519 1538 -3850 1558
rect -6519 1536 -4060 1538
rect -6309 1481 -4060 1536
rect -6309 1479 -3850 1481
rect -6519 1469 -3850 1479
rect -9457 1421 -9447 1439
rect -10115 824 -9447 1421
rect -10115 640 -10109 824
rect -9457 640 -9447 824
rect -9395 640 -9385 1439
rect -8687 1398 -6519 1404
rect -8689 1392 -6519 1398
rect -6309 1398 -6299 1404
rect -6229 1398 -6219 1403
rect -8689 1358 -8677 1392
rect -8689 1352 -6519 1358
rect -8687 1347 -6519 1352
rect -6309 1352 -6297 1398
rect -6231 1352 -6219 1398
rect -6009 1398 -3841 1403
rect -6009 1392 -3839 1398
rect -3851 1358 -3839 1392
rect -6309 1347 -6299 1352
rect -8745 1308 -8699 1320
rect -10155 628 -10109 640
rect -9445 628 -9386 640
rect -10077 612 -9477 618
rect -10077 578 -10065 612
rect -9489 578 -9477 612
rect -10077 572 -9477 578
rect -8898 236 -8849 1308
rect -8697 236 -8687 1308
rect -8898 167 -8739 236
rect -8745 132 -8739 167
rect -8705 167 -8687 236
rect -8705 132 -8699 167
rect -8745 120 -8699 132
rect -8045 89 -6958 1347
rect -6229 1346 -6219 1352
rect -6009 1352 -3839 1358
rect -6009 1346 -3841 1352
rect -6287 1308 -6241 1320
rect -6287 1277 -6281 1308
rect -6247 1277 -6241 1308
rect -6299 958 -6289 1277
rect -6237 958 -6227 1277
rect -6287 132 -6281 958
rect -6247 132 -6241 958
rect -6287 120 -6241 132
rect -10303 68 -9726 74
rect -10303 -26 -10291 68
rect -9738 -26 -9726 68
rect -8689 37 -8677 89
rect -8197 82 -6297 89
rect -6229 88 -6219 90
rect -6309 48 -6297 82
rect -8197 37 -6297 48
rect -6231 42 -6219 88
rect -5739 88 -5729 90
rect -5545 88 -4458 1346
rect -3829 1308 -3783 1320
rect -3842 236 -3832 1308
rect -3680 236 -3670 1308
rect -3829 132 -3823 236
rect -3789 132 -3783 236
rect -3829 120 -3783 132
rect -5739 82 -3839 88
rect -3851 48 -3839 82
rect -6229 38 -6219 42
rect -5739 42 -3839 48
rect -5739 38 -5729 42
rect -1807 22 -1797 3198
rect -10303 -32 -9726 -26
rect -1808 -154 -1798 22
rect -1649 -5 -1639 3198
rect -1482 3154 -1436 3166
rect -1501 2154 -1491 3154
rect -1427 2154 -1417 3154
rect -1482 178 -1476 2154
rect -1442 178 -1436 2154
rect -1482 166 -1436 178
rect -1350 125 -1145 3204
rect -1044 3154 -998 3166
rect -1044 778 -1038 3154
rect -1004 778 -998 3154
rect -1067 178 -1057 778
rect -985 178 -975 778
rect -1044 166 -998 178
rect -897 125 -692 3204
rect -606 3154 -560 3166
rect -606 1994 -600 3154
rect -566 1994 -560 3154
rect -625 994 -615 1994
rect -551 994 -541 1994
rect -606 178 -600 994
rect -566 178 -560 994
rect -606 166 -560 178
rect -461 125 -256 3204
rect -168 3154 -122 3166
rect -168 778 -162 3154
rect -128 778 -122 3154
rect -192 178 -182 778
rect -110 178 -100 778
rect -168 166 -122 178
rect -29 125 176 3204
rect 270 3154 316 3166
rect 251 2154 261 3154
rect 325 2154 335 3154
rect 11783 2778 12054 2785
rect 7074 2773 12054 2778
rect 7074 2772 11789 2773
rect 576 2612 730 2624
rect 270 178 276 2154
rect 310 178 316 2154
rect 270 166 316 178
rect 576 132 582 2612
rect 724 2120 730 2612
rect 7074 2407 7086 2772
rect 12048 2408 12058 2773
rect 11890 2407 11932 2408
rect 7074 2401 7148 2407
rect 5231 2120 5530 2125
rect 724 2114 5530 2120
rect 5514 2113 5530 2114
rect 724 1816 2986 1822
rect 724 132 730 1816
rect -1426 119 -1054 125
rect -1426 85 -1414 119
rect -1066 85 -1054 119
rect -1426 79 -1054 85
rect -988 119 -616 125
rect -988 85 -976 119
rect -628 85 -616 119
rect -988 79 -616 85
rect -550 119 -178 125
rect -550 85 -538 119
rect -190 85 -178 119
rect -550 79 -178 85
rect -112 119 260 125
rect 576 120 730 132
rect -112 85 -100 119
rect 248 85 260 119
rect -112 79 260 85
rect -1649 -11 779 -5
rect -1804 -155 -1685 -154
rect 767 -155 779 -11
rect -1804 -161 779 -155
rect -10301 -167 -3343 -161
rect -1804 -166 -1643 -161
rect -10301 -256 -10289 -167
rect -3355 -256 -3343 -167
rect 2980 -168 2986 1816
rect 3219 1816 5237 1822
rect 3219 72 3225 1816
rect 3403 1693 3755 1699
rect 3403 1659 3415 1693
rect 3743 1659 3755 1693
rect 3403 1653 3755 1659
rect 3821 1693 4173 1699
rect 3821 1659 3833 1693
rect 4161 1659 4173 1693
rect 3821 1653 4173 1659
rect 4239 1693 4591 1699
rect 4239 1659 4251 1693
rect 4579 1659 4591 1693
rect 4239 1653 4591 1659
rect 4657 1693 5009 1699
rect 4657 1659 4669 1693
rect 4997 1659 5009 1693
rect 4657 1653 5009 1659
rect 3347 1600 3393 1612
rect 3334 600 3344 1600
rect 3396 600 3406 1600
rect 3347 224 3353 600
rect 3387 224 3393 600
rect 3347 212 3393 224
rect 3471 171 3672 1653
rect 3765 1600 3811 1612
rect 3765 1224 3771 1600
rect 3805 1224 3811 1600
rect 3752 224 3762 1224
rect 3814 224 3824 1224
rect 3765 212 3811 224
rect 3890 171 4091 1653
rect 4183 1600 4229 1612
rect 4170 600 4180 1600
rect 4232 600 4242 1600
rect 4183 224 4189 600
rect 4223 224 4229 600
rect 4183 212 4229 224
rect 4313 171 4514 1653
rect 4601 1600 4647 1612
rect 4601 1224 4607 1600
rect 4641 1224 4647 1600
rect 4588 224 4598 1224
rect 4650 224 4660 1224
rect 4601 212 4647 224
rect 4719 171 4920 1653
rect 5019 1600 5065 1612
rect 5006 600 5016 1600
rect 5068 600 5078 1600
rect 5019 224 5025 600
rect 5059 224 5065 600
rect 5227 306 5237 1816
rect 5524 306 5534 2113
rect 5231 294 5530 306
rect 5019 212 5065 224
rect 5214 171 5224 180
rect 3403 165 5224 171
rect 3403 131 3415 165
rect 3743 131 3833 165
rect 4161 131 4251 165
rect 4579 131 4669 165
rect 4997 131 5224 165
rect 3403 125 5224 131
rect 5214 121 5224 125
rect 5348 121 5358 180
rect 7138 115 7148 2401
rect 7265 2401 11932 2407
rect 7265 211 7275 2401
rect 11783 2396 11932 2401
rect 7440 2238 8488 2244
rect 7440 2204 7508 2238
rect 8476 2204 8488 2238
rect 7440 2198 8488 2204
rect 8554 2238 10604 2244
rect 8554 2204 8566 2238
rect 9534 2204 9624 2238
rect 10592 2204 10604 2238
rect 8554 2198 10604 2204
rect 10670 2238 11718 2244
rect 10670 2204 10682 2238
rect 11650 2204 11718 2238
rect 10670 2198 11718 2204
rect 7440 2145 7486 2198
rect 8498 2145 8544 2157
rect 9556 2145 9602 2198
rect 10614 2145 10660 2157
rect 11672 2145 11718 2198
rect 7440 1869 7446 2145
rect 7480 1869 7486 2145
rect 7421 1669 7431 1869
rect 7495 1669 7505 1869
rect 8485 1845 8495 2145
rect 8547 1845 8557 2145
rect 9537 1945 9547 2145
rect 9611 1945 9621 2145
rect 8498 1669 8504 1845
rect 8538 1669 8544 1845
rect 7440 1616 7486 1669
rect 8498 1657 8544 1669
rect 9556 1669 9562 1945
rect 9596 1669 9602 1945
rect 10601 1845 10611 2145
rect 10663 1845 10673 2145
rect 11672 1869 11678 2145
rect 11712 1869 11718 2145
rect 9556 1619 9602 1669
rect 10614 1669 10620 1845
rect 10654 1669 10660 1845
rect 11653 1669 11663 1869
rect 11727 1669 11737 1869
rect 10614 1657 10660 1669
rect 11672 1657 11718 1669
rect 7826 1616 7836 1619
rect 7440 1610 7836 1616
rect 8476 1616 8486 1619
rect 8884 1616 8894 1619
rect 7440 1576 7508 1610
rect 7440 1570 7836 1576
rect 7826 1567 7836 1570
rect 8476 1570 8488 1616
rect 8554 1610 8894 1616
rect 9534 1616 9617 1619
rect 9942 1616 9952 1620
rect 9534 1610 9952 1616
rect 10592 1616 10602 1620
rect 11000 1616 11010 1619
rect 8554 1576 8566 1610
rect 9534 1576 9624 1610
rect 8554 1570 8894 1576
rect 8476 1567 8486 1570
rect 8884 1567 8894 1570
rect 9534 1570 9952 1576
rect 9534 1567 9617 1570
rect 9942 1568 9952 1570
rect 10592 1570 10604 1616
rect 10670 1610 11010 1616
rect 11650 1616 11660 1619
rect 10670 1576 10682 1610
rect 10670 1570 11010 1576
rect 10592 1568 10602 1570
rect 11000 1567 11010 1570
rect 11650 1570 11662 1616
rect 11922 1594 11932 2396
rect 12029 2396 12054 2408
rect 12029 1594 12039 2396
rect 11926 1582 12035 1594
rect 11650 1567 11660 1570
rect 7489 1371 8376 1471
rect 8476 1371 8566 1471
rect 8666 1371 9624 1471
rect 9724 1371 11550 1471
rect 11650 1371 12265 1471
rect 7492 1189 7508 1289
rect 7608 1189 9434 1289
rect 9534 1189 10492 1289
rect 10592 1189 10682 1289
rect 10782 1189 11910 1289
rect 7440 1085 7486 1086
rect 7440 1033 7508 1085
rect 8148 1082 8158 1085
rect 8556 1082 8566 1085
rect 8148 1076 8488 1082
rect 8476 1042 8488 1076
rect 8148 1036 8488 1042
rect 8554 1036 8566 1082
rect 9206 1082 9216 1085
rect 9614 1082 9624 1085
rect 9206 1076 9624 1082
rect 10264 1082 10274 1085
rect 10672 1082 10682 1085
rect 10264 1076 10604 1082
rect 9534 1042 9624 1076
rect 10592 1042 10604 1076
rect 8148 1033 8158 1036
rect 8556 1033 8566 1036
rect 9206 1036 9624 1042
rect 9206 1033 9216 1036
rect 9556 1033 9624 1036
rect 10264 1036 10604 1042
rect 10670 1036 10682 1082
rect 11322 1082 11332 1085
rect 11322 1076 11718 1082
rect 11650 1042 11718 1076
rect 10264 1033 10274 1036
rect 10672 1033 10682 1036
rect 11322 1036 11718 1042
rect 11322 1033 11332 1036
rect 7440 1032 7518 1033
rect 7440 983 7486 1032
rect 8498 983 8544 995
rect 7421 783 7431 983
rect 7495 783 7505 983
rect 8498 807 8504 983
rect 8538 807 8544 983
rect 9556 983 9602 1033
rect 7440 507 7446 783
rect 7480 507 7486 783
rect 8485 507 8495 807
rect 8547 507 8557 807
rect 9556 707 9562 983
rect 9596 707 9602 983
rect 10614 983 10660 995
rect 11672 983 11718 1036
rect 10614 807 10620 983
rect 10654 807 10660 983
rect 9537 507 9547 707
rect 9611 507 9621 707
rect 10601 507 10611 807
rect 10663 507 10673 807
rect 11653 783 11663 983
rect 11727 783 11737 983
rect 11672 507 11678 783
rect 11712 507 11718 783
rect 7440 454 7486 507
rect 8498 495 8544 507
rect 9556 454 9602 507
rect 10614 495 10660 507
rect 11672 454 11718 507
rect 7440 448 8488 454
rect 7440 414 7508 448
rect 8476 414 8488 448
rect 7440 408 8488 414
rect 8554 448 10604 454
rect 8554 414 8566 448
rect 9534 414 9624 448
rect 10592 414 10604 448
rect 8554 408 10604 414
rect 10670 448 11718 454
rect 10670 414 10682 448
rect 11650 414 11718 448
rect 10670 408 11718 414
rect 7265 205 11709 211
rect 7142 108 7183 115
rect 7142 103 11593 108
rect 7171 102 11593 103
rect 3219 66 5146 72
rect 2980 -170 3071 -168
rect 5134 -170 5146 66
rect 8500 -19 8570 -13
rect 10573 -19 10661 -13
rect 8500 -25 10661 -19
rect 2980 -176 5146 -170
rect 2980 -180 3225 -176
rect -10301 -262 -3343 -256
rect 6078 -456 6206 -437
rect -1748 -493 -1589 -481
rect -1752 -1789 -1742 -493
rect -1595 -495 -1585 -493
rect -1595 -496 -1454 -495
rect 6068 -496 6078 -456
rect -1595 -501 6078 -496
rect -1466 -502 6078 -501
rect -1754 -1993 -1742 -1789
rect -1595 -611 6078 -605
rect -1595 -1789 -1585 -611
rect 6068 -639 6078 -611
rect 6225 -639 6235 -456
rect 8496 -666 8506 -25
rect 8564 -134 10579 -128
rect 8564 -666 8574 -134
rect 8681 -218 9073 -212
rect 8681 -252 8693 -218
rect 9061 -252 9073 -218
rect 8681 -258 9073 -252
rect 9139 -218 9531 -212
rect 9139 -252 9151 -218
rect 9519 -252 9531 -218
rect 9139 -258 9531 -252
rect 9597 -218 9989 -212
rect 9597 -252 9609 -218
rect 9977 -252 9989 -218
rect 9597 -258 9989 -252
rect 10055 -218 10447 -212
rect 10055 -252 10067 -218
rect 10435 -252 10447 -218
rect 10055 -258 10447 -252
rect 8625 -302 8671 -290
rect 9083 -302 9129 -290
rect 9541 -302 9587 -290
rect 9999 -302 10045 -290
rect 10457 -302 10503 -290
rect 8500 -678 8570 -666
rect 8625 -731 8631 -302
rect 8665 -731 8671 -302
rect 9070 -462 9080 -302
rect 9132 -462 9142 -302
rect -1416 -788 456 -782
rect -1416 -822 -1404 -788
rect 444 -822 456 -788
rect -1416 -828 456 -822
rect 522 -788 4332 -782
rect 522 -822 534 -788
rect 2382 -822 2472 -788
rect 4320 -822 4332 -788
rect 522 -828 4332 -822
rect 4398 -788 6270 -782
rect 4398 -822 4410 -788
rect 6258 -822 6270 -788
rect 4398 -828 6270 -822
rect -1472 -872 -1426 -860
rect -1491 -972 -1481 -872
rect -1417 -972 -1407 -872
rect -1472 -1148 -1466 -972
rect -1432 -1148 -1426 -972
rect -1472 -1160 -1426 -1148
rect -1196 -1192 223 -828
rect 466 -872 512 -860
rect 453 -972 463 -872
rect 515 -972 525 -872
rect 466 -1148 472 -972
rect 506 -1148 512 -972
rect 466 -1160 512 -1148
rect 838 -1192 2257 -828
rect 2404 -872 2450 -828
rect 2404 -1048 2410 -872
rect 2444 -1048 2450 -872
rect 2385 -1148 2395 -1048
rect 2459 -1148 2469 -1048
rect 2404 -1160 2450 -1148
rect 2667 -1192 4086 -828
rect 4342 -872 4388 -860
rect 4329 -972 4339 -872
rect 4391 -972 4401 -872
rect 4342 -1148 4348 -972
rect 4382 -1148 4388 -972
rect 4342 -1160 4388 -1148
rect 4637 -1192 6056 -828
rect 6280 -872 6326 -860
rect 8589 -868 8599 -731
rect 8693 -868 8703 -731
rect 6261 -972 6271 -872
rect 6335 -972 6345 -872
rect 8625 -878 8631 -868
rect 8665 -878 8671 -868
rect 8625 -890 8671 -878
rect 9083 -878 9089 -462
rect 9123 -878 9129 -462
rect 9541 -473 9547 -302
rect 9581 -473 9587 -302
rect 9986 -462 9996 -302
rect 10048 -462 10058 -302
rect 9508 -610 9518 -473
rect 9612 -610 9622 -473
rect 9083 -890 9129 -878
rect 9541 -878 9547 -610
rect 9581 -878 9587 -610
rect 9541 -890 9587 -878
rect 9999 -878 10005 -462
rect 10039 -878 10045 -462
rect 10457 -731 10463 -302
rect 10497 -731 10503 -302
rect 10424 -868 10434 -731
rect 10528 -868 10538 -731
rect 9999 -890 10045 -878
rect 10457 -878 10463 -868
rect 10497 -878 10503 -868
rect 10457 -890 10503 -878
rect 8851 -922 8861 -919
rect 8681 -928 8861 -922
rect 9061 -922 9071 -919
rect 9309 -922 9319 -919
rect 8681 -962 8693 -928
rect 8681 -968 8861 -962
rect 8851 -971 8861 -968
rect 9061 -968 9073 -922
rect 9139 -928 9319 -922
rect 9519 -922 9529 -919
rect 9767 -922 9777 -919
rect 9139 -962 9151 -928
rect 9139 -968 9319 -962
rect 9061 -971 9071 -968
rect 9309 -971 9319 -968
rect 9519 -968 9531 -922
rect 9597 -928 9777 -922
rect 9977 -922 9987 -919
rect 10225 -922 10235 -919
rect 9597 -962 9609 -928
rect 9597 -968 9777 -962
rect 9519 -971 9529 -968
rect 9767 -971 9777 -968
rect 9977 -968 9989 -922
rect 10055 -928 10235 -922
rect 10435 -922 10445 -919
rect 10055 -962 10067 -928
rect 10055 -968 10235 -962
rect 9977 -971 9987 -968
rect 10225 -971 10235 -968
rect 10435 -968 10447 -922
rect 10435 -971 10445 -968
rect 6280 -1148 6286 -972
rect 6320 -1148 6326 -972
rect 7112 -1143 7122 -1043
rect 7205 -1143 8961 -1043
rect 9061 -1143 9151 -1043
rect 9251 -1143 9609 -1043
rect 9709 -1143 10335 -1043
rect 10435 -1143 10480 -1043
rect 6280 -1160 6326 -1148
rect -1416 -1198 6270 -1192
rect -1416 -1232 -1404 -1198
rect 444 -1232 534 -1198
rect 2382 -1232 2472 -1198
rect 4320 -1232 4410 -1198
rect 6258 -1232 6270 -1198
rect -1416 -1238 6270 -1232
rect -1472 -1282 -1426 -1270
rect -1472 -1458 -1466 -1282
rect -1432 -1458 -1426 -1282
rect -1491 -1558 -1481 -1458
rect -1417 -1558 -1407 -1458
rect -1472 -1602 -1426 -1558
rect -1192 -1602 227 -1238
rect 466 -1282 512 -1270
rect 466 -1458 472 -1282
rect 506 -1458 512 -1282
rect 453 -1558 463 -1458
rect 515 -1558 525 -1458
rect 466 -1570 512 -1558
rect 834 -1602 2253 -1238
rect 2404 -1282 2450 -1270
rect 2385 -1382 2395 -1282
rect 2459 -1382 2469 -1282
rect 2404 -1558 2410 -1382
rect 2444 -1558 2450 -1382
rect 2404 -1570 2450 -1558
rect 2667 -1602 4086 -1238
rect 4342 -1282 4388 -1270
rect 4342 -1458 4348 -1282
rect 4382 -1458 4388 -1282
rect 4329 -1558 4339 -1458
rect 4391 -1558 4401 -1458
rect 4342 -1570 4388 -1558
rect 4637 -1602 6056 -1238
rect 6280 -1282 6326 -1270
rect 6280 -1458 6286 -1282
rect 6320 -1458 6326 -1282
rect 7102 -1329 7112 -1229
rect 7225 -1329 8693 -1229
rect 8793 -1329 9419 -1229
rect 9519 -1329 9877 -1229
rect 9977 -1329 10067 -1229
rect 10167 -1329 10480 -1229
rect 8683 -1419 8693 -1416
rect 6261 -1558 6271 -1458
rect 6335 -1558 6345 -1458
rect 8681 -1465 8693 -1419
rect 8893 -1419 8903 -1416
rect 9141 -1419 9151 -1416
rect 8893 -1425 9073 -1419
rect 9061 -1459 9073 -1425
rect 8683 -1468 8693 -1465
rect 8893 -1465 9073 -1459
rect 9139 -1465 9151 -1419
rect 9351 -1419 9361 -1416
rect 9599 -1419 9609 -1416
rect 9351 -1425 9531 -1419
rect 9519 -1459 9531 -1425
rect 8893 -1468 8903 -1465
rect 9141 -1468 9151 -1465
rect 9351 -1465 9531 -1459
rect 9597 -1465 9609 -1419
rect 9809 -1419 9819 -1416
rect 10057 -1419 10067 -1416
rect 9809 -1425 9989 -1419
rect 9977 -1459 9989 -1425
rect 9351 -1468 9361 -1465
rect 9599 -1468 9609 -1465
rect 9809 -1465 9989 -1459
rect 10055 -1465 10067 -1419
rect 10267 -1419 10277 -1416
rect 10267 -1425 10447 -1419
rect 10435 -1459 10447 -1425
rect 9809 -1468 9819 -1465
rect 10057 -1468 10067 -1465
rect 10267 -1465 10447 -1459
rect 10267 -1468 10277 -1465
rect 8625 -1509 8671 -1497
rect 8625 -1520 8631 -1509
rect 8665 -1520 8671 -1509
rect 9083 -1509 9129 -1497
rect 6280 -1602 6326 -1558
rect -1472 -1608 456 -1602
rect -1472 -1642 -1404 -1608
rect 444 -1642 456 -1608
rect -1472 -1648 456 -1642
rect 522 -1608 2394 -1602
rect 522 -1642 534 -1608
rect 2382 -1642 2394 -1608
rect 522 -1648 2394 -1642
rect 2460 -1608 4332 -1602
rect 2460 -1642 2472 -1608
rect 4320 -1642 4332 -1608
rect 2460 -1648 4332 -1642
rect 4398 -1608 6326 -1602
rect 4398 -1642 4410 -1608
rect 6258 -1642 6326 -1608
rect 4398 -1648 6326 -1642
rect 8590 -1657 8600 -1520
rect 8694 -1657 8704 -1520
rect 8491 -1702 8577 -1690
rect -1595 -1790 -1489 -1789
rect -1595 -1795 6189 -1790
rect -1501 -1796 6189 -1795
rect 6177 -1993 6189 -1796
rect -1754 -1999 6189 -1993
rect 8487 -2321 8497 -1702
rect 8446 -2333 8497 -2321
rect 8571 -2321 8581 -1702
rect 8625 -2085 8631 -1657
rect 8665 -2085 8671 -1657
rect 9083 -1925 9089 -1509
rect 9123 -1925 9129 -1509
rect 9541 -1509 9587 -1497
rect 9541 -1731 9547 -1509
rect 9581 -1731 9587 -1509
rect 9999 -1509 10045 -1497
rect 9507 -1868 9517 -1731
rect 9611 -1868 9621 -1731
rect 9070 -2085 9080 -1925
rect 9132 -2085 9142 -1925
rect 9541 -2085 9547 -1868
rect 9581 -2085 9587 -1868
rect 9999 -1925 10005 -1509
rect 10039 -1925 10045 -1509
rect 10457 -1509 10503 -1497
rect 10457 -1520 10463 -1509
rect 10497 -1520 10503 -1509
rect 10422 -1657 10432 -1520
rect 10526 -1657 10536 -1520
rect 9986 -2085 9996 -1925
rect 10048 -2085 10058 -1925
rect 10457 -2085 10463 -1657
rect 10497 -2085 10503 -1657
rect 8625 -2097 8671 -2085
rect 9083 -2097 9129 -2085
rect 9541 -2097 9587 -2085
rect 9999 -2097 10045 -2085
rect 10457 -2097 10503 -2085
rect 8681 -2135 9073 -2129
rect 8681 -2169 8693 -2135
rect 9061 -2169 9073 -2135
rect 8681 -2175 9073 -2169
rect 9139 -2135 9531 -2129
rect 9139 -2169 9151 -2135
rect 9519 -2169 9531 -2135
rect 9139 -2175 9531 -2169
rect 9597 -2135 9989 -2129
rect 9597 -2169 9609 -2135
rect 9977 -2169 9989 -2135
rect 9597 -2175 9989 -2169
rect 10055 -2135 10447 -2129
rect 10055 -2169 10067 -2135
rect 10435 -2169 10447 -2135
rect 10055 -2175 10447 -2169
rect 8571 -2327 8685 -2321
rect 10573 -2327 10579 -134
rect 8571 -2333 10579 -2327
rect 10655 -2327 10661 -25
rect 11583 -1051 11593 102
rect 11697 102 11709 205
rect 11697 -1051 11707 102
rect 11810 -327 11910 1189
rect 11810 -361 11841 -327
rect 11879 -361 11910 -327
rect 11810 -367 11910 -361
rect 12165 -327 12265 1371
rect 12165 -361 12197 -327
rect 12235 -361 12265 -327
rect 12165 -367 12265 -361
rect 11773 -420 11819 -408
rect 11901 -420 11947 -408
rect 12129 -420 12175 -408
rect 12257 -420 12303 -408
rect 11760 -620 11770 -420
rect 11822 -620 11832 -420
rect 11773 -916 11779 -620
rect 11813 -916 11819 -620
rect 11901 -716 11907 -420
rect 11941 -716 11947 -420
rect 12116 -620 12126 -420
rect 12178 -620 12188 -420
rect 11888 -916 11898 -716
rect 11950 -916 11960 -716
rect 12129 -916 12135 -620
rect 12169 -916 12175 -620
rect 12257 -716 12263 -420
rect 12297 -716 12303 -420
rect 12244 -916 12254 -716
rect 12306 -916 12316 -716
rect 11773 -928 11819 -916
rect 11901 -928 11947 -916
rect 12129 -928 12175 -916
rect 12257 -928 12303 -916
rect 11827 -975 11892 -968
rect 11827 -1009 11841 -975
rect 11879 -1009 11892 -975
rect 11827 -1026 11892 -1009
rect 12185 -975 12247 -969
rect 12185 -1009 12197 -975
rect 12235 -1009 12247 -975
rect 12185 -1040 12247 -1009
rect 11587 -1063 11703 -1051
rect 11888 -1335 11898 -1302
rect 11851 -1341 11898 -1335
rect 11851 -1375 11863 -1341
rect 11897 -1375 11898 -1341
rect 11851 -1381 11898 -1375
rect 11950 -1335 11960 -1302
rect 11950 -1341 12265 -1335
rect 11950 -1375 12219 -1341
rect 12253 -1375 12265 -1341
rect 11950 -1381 12265 -1375
rect 11907 -1413 11941 -1381
rect 11813 -1425 11859 -1413
rect 11813 -1530 11819 -1425
rect 11853 -1530 11859 -1425
rect 11901 -1425 11947 -1413
rect 11800 -1601 11810 -1530
rect 11862 -1601 11872 -1530
rect 11901 -1601 11907 -1425
rect 11941 -1601 11947 -1425
rect 12169 -1425 12215 -1413
rect 12257 -1425 12303 -1413
rect 12169 -1530 12175 -1425
rect 12209 -1530 12215 -1425
rect 12244 -1496 12254 -1425
rect 12306 -1496 12316 -1425
rect 12156 -1601 12166 -1530
rect 12218 -1601 12228 -1530
rect 12257 -1601 12263 -1496
rect 12297 -1601 12303 -1496
rect 11813 -1613 11859 -1601
rect 11901 -1613 11947 -1601
rect 12169 -1613 12215 -1601
rect 12257 -1613 12303 -1601
rect 11851 -1651 12265 -1645
rect 11851 -1685 11863 -1651
rect 11897 -1685 12219 -1651
rect 12253 -1685 12265 -1651
rect 11851 -1691 12265 -1685
rect 10985 -1885 12387 -1879
rect 10985 -2163 10997 -1885
rect 12375 -2157 12387 -1885
rect 10991 -2321 10997 -2163
rect 10922 -2327 10997 -2321
rect 10655 -2333 10997 -2327
rect 11117 -2163 12387 -2157
rect 3710 -2888 3861 -2878
rect 2116 -2918 2319 -2906
rect -1567 -3685 -1381 -3673
rect -1567 -10263 -1561 -3685
rect -1387 -10263 -1381 -3685
rect 1374 -3729 1498 -3717
rect -1136 -3800 -936 -3790
rect -1148 -3855 -1136 -3809
rect 921 -3806 1121 -3796
rect -936 -3815 -348 -3809
rect -360 -3849 -348 -3815
rect 333 -3815 921 -3809
rect -936 -3855 -348 -3849
rect -93 -3829 -41 -3819
rect -1226 -3877 -1180 -3865
rect -1136 -3874 -936 -3864
rect -316 -3867 -270 -3865
rect -1226 -4045 -1220 -3877
rect -1186 -3916 -1180 -3877
rect -319 -3877 -267 -3867
rect -1186 -3977 -319 -3916
rect -1186 -4004 -310 -3977
rect -1186 -4045 -1180 -4004
rect -1226 -4135 -1180 -4045
rect -316 -4045 -310 -4004
rect -276 -3987 -267 -3977
rect -276 -4045 -270 -3987
rect -560 -4062 -360 -4052
rect -1148 -4073 -560 -4067
rect -1148 -4107 -1136 -4073
rect -1148 -4113 -560 -4107
rect -360 -4113 -348 -4067
rect -560 -4128 -360 -4118
rect -1226 -4303 -1220 -4135
rect -1186 -4159 -1180 -4135
rect -316 -4135 -270 -4045
rect -316 -4159 -310 -4135
rect -1186 -4247 -310 -4159
rect -1186 -4303 -1180 -4247
rect -1226 -4315 -1180 -4303
rect -316 -4303 -310 -4247
rect -276 -4303 -270 -4135
rect -784 -4322 -684 -4312
rect -316 -4315 -270 -4303
rect -93 -4087 -41 -3929
rect -1148 -4331 -784 -4325
rect -684 -4331 -348 -4325
rect -1148 -4365 -1136 -4331
rect -360 -4365 -348 -4331
rect -1148 -4371 -784 -4365
rect -684 -4371 -348 -4365
rect -1226 -4393 -1180 -4381
rect -784 -4384 -684 -4374
rect -316 -4383 -270 -4381
rect -1226 -4561 -1220 -4393
rect -1186 -4433 -1180 -4393
rect -319 -4393 -267 -4383
rect -1186 -4451 -319 -4433
rect -1186 -4503 -790 -4451
rect -685 -4493 -319 -4451
rect -685 -4503 -310 -4493
rect -1186 -4521 -310 -4503
rect -1186 -4561 -1180 -4521
rect -1226 -4651 -1180 -4561
rect -316 -4561 -310 -4521
rect -276 -4503 -267 -4493
rect -276 -4561 -270 -4503
rect -1136 -4580 -936 -4570
rect -1148 -4629 -1136 -4583
rect -936 -4589 -348 -4583
rect -360 -4623 -348 -4589
rect -936 -4629 -348 -4623
rect -1136 -4642 -936 -4632
rect -1226 -4819 -1220 -4651
rect -1186 -4690 -1180 -4651
rect -316 -4651 -270 -4561
rect -316 -4690 -310 -4651
rect -1186 -4713 -310 -4690
rect -1186 -4765 -787 -4713
rect -687 -4765 -310 -4713
rect -1186 -4778 -310 -4765
rect -1186 -4819 -1180 -4778
rect -1226 -4831 -1180 -4819
rect -316 -4819 -310 -4778
rect -276 -4819 -270 -4651
rect -784 -4838 -684 -4828
rect -316 -4831 -270 -4819
rect -1148 -4847 -784 -4841
rect -684 -4847 -348 -4841
rect -1148 -4881 -1136 -4847
rect -360 -4881 -348 -4847
rect -1148 -4887 -784 -4881
rect -684 -4887 -348 -4881
rect -93 -4861 -41 -4187
rect -1226 -4909 -1180 -4897
rect -784 -4900 -684 -4890
rect -316 -4899 -270 -4897
rect -1226 -5077 -1220 -4909
rect -1186 -4956 -1180 -4909
rect -319 -4909 -267 -4899
rect -1186 -5034 -319 -4956
rect -1186 -5044 -310 -5034
rect -1186 -5077 -1180 -5044
rect -1226 -5167 -1180 -5077
rect -316 -5077 -310 -5044
rect -276 -5040 -267 -5034
rect -276 -5077 -270 -5040
rect -560 -5094 -360 -5084
rect -1148 -5105 -560 -5099
rect -1148 -5139 -1136 -5105
rect -1148 -5145 -560 -5139
rect -360 -5145 -348 -5099
rect -560 -5160 -360 -5150
rect -1226 -5335 -1220 -5167
rect -1186 -5207 -1180 -5167
rect -316 -5167 -270 -5077
rect -316 -5207 -310 -5167
rect -1186 -5295 -310 -5207
rect -1186 -5335 -1180 -5295
rect -1226 -5425 -1180 -5335
rect -316 -5335 -310 -5295
rect -276 -5335 -270 -5167
rect -1136 -5348 -936 -5338
rect -1148 -5403 -1136 -5357
rect -936 -5363 -348 -5357
rect -360 -5397 -348 -5363
rect -936 -5403 -348 -5397
rect -1136 -5422 -936 -5412
rect -1226 -5593 -1220 -5425
rect -1186 -5472 -1180 -5425
rect -316 -5425 -270 -5335
rect -316 -5472 -310 -5425
rect -1186 -5560 -310 -5472
rect -1186 -5593 -1180 -5560
rect -1226 -5683 -1180 -5593
rect -316 -5593 -310 -5560
rect -276 -5593 -270 -5425
rect -560 -5610 -360 -5600
rect -1148 -5621 -560 -5615
rect -1148 -5655 -1136 -5621
rect -1148 -5661 -560 -5655
rect -360 -5661 -348 -5615
rect -560 -5676 -360 -5666
rect -1226 -5851 -1220 -5683
rect -1186 -5716 -1180 -5683
rect -316 -5683 -270 -5593
rect -316 -5716 -310 -5683
rect -1186 -5804 -310 -5716
rect -1186 -5851 -1180 -5804
rect -1226 -5863 -1180 -5851
rect -316 -5851 -310 -5804
rect -276 -5851 -270 -5683
rect -784 -5870 -684 -5860
rect -316 -5863 -270 -5851
rect -93 -5635 -41 -4961
rect -1148 -5879 -784 -5873
rect -684 -5879 -348 -5873
rect -1148 -5913 -1136 -5879
rect -360 -5913 -348 -5879
rect -1148 -5919 -784 -5913
rect -684 -5919 -348 -5913
rect -1226 -5941 -1180 -5929
rect -784 -5932 -684 -5922
rect -316 -5931 -270 -5929
rect -1226 -6109 -1220 -5941
rect -1186 -5983 -1180 -5941
rect -319 -5941 -267 -5931
rect -1186 -6004 -319 -5983
rect -1186 -6056 -785 -6004
rect -685 -6041 -319 -6004
rect -685 -6056 -310 -6041
rect -1186 -6071 -310 -6056
rect -1186 -6109 -1180 -6071
rect -1226 -6199 -1180 -6109
rect -316 -6109 -310 -6071
rect -276 -6051 -267 -6041
rect -276 -6109 -270 -6051
rect -1136 -6129 -936 -6119
rect -1148 -6177 -1136 -6131
rect -936 -6137 -348 -6131
rect -360 -6171 -348 -6137
rect -936 -6177 -348 -6171
rect -1136 -6191 -936 -6181
rect -1226 -6367 -1220 -6199
rect -1186 -6240 -1180 -6199
rect -316 -6199 -270 -6109
rect -316 -6240 -310 -6199
rect -1186 -6256 -310 -6240
rect -1186 -6308 -782 -6256
rect -682 -6308 -310 -6256
rect -1186 -6328 -310 -6308
rect -1186 -6367 -1180 -6328
rect -1226 -6379 -1180 -6367
rect -316 -6367 -310 -6328
rect -276 -6367 -270 -6199
rect -784 -6386 -684 -6376
rect -316 -6379 -270 -6367
rect -1148 -6395 -784 -6389
rect -684 -6395 -348 -6389
rect -1148 -6429 -1136 -6395
rect -360 -6429 -348 -6395
rect -1148 -6435 -784 -6429
rect -684 -6435 -348 -6429
rect -93 -6409 -41 -5735
rect -1226 -6457 -1180 -6445
rect -784 -6448 -684 -6438
rect -316 -6447 -270 -6445
rect -1226 -6625 -1220 -6457
rect -1186 -6492 -1180 -6457
rect -319 -6457 -267 -6447
rect -1186 -6580 -319 -6492
rect -1186 -6625 -1180 -6580
rect -319 -6597 -310 -6583
rect -1226 -6715 -1180 -6625
rect -316 -6625 -310 -6597
rect -276 -6597 -267 -6583
rect -276 -6625 -270 -6597
rect -560 -6642 -360 -6632
rect -1148 -6653 -560 -6647
rect -1148 -6687 -1136 -6653
rect -1148 -6693 -560 -6687
rect -360 -6693 -348 -6647
rect -560 -6708 -360 -6698
rect -1226 -6883 -1220 -6715
rect -1186 -6751 -1180 -6715
rect -316 -6715 -270 -6625
rect -316 -6751 -310 -6715
rect -1186 -6839 -310 -6751
rect -1186 -6883 -1180 -6839
rect -1226 -6973 -1180 -6883
rect -316 -6883 -310 -6839
rect -276 -6883 -270 -6715
rect -1136 -6896 -936 -6886
rect -1148 -6951 -1136 -6905
rect -936 -6911 -348 -6905
rect -360 -6945 -348 -6911
rect -936 -6951 -348 -6945
rect -1136 -6970 -936 -6960
rect -1226 -7141 -1220 -6973
rect -1186 -7008 -1180 -6973
rect -316 -6973 -270 -6883
rect -316 -7008 -310 -6973
rect -1186 -7096 -310 -7008
rect -1186 -7141 -1180 -7096
rect -1226 -7231 -1180 -7141
rect -316 -7141 -310 -7096
rect -276 -7141 -270 -6973
rect -560 -7158 -360 -7148
rect -1148 -7169 -560 -7163
rect -1148 -7203 -1136 -7169
rect -1148 -7209 -560 -7203
rect -360 -7209 -348 -7163
rect -560 -7224 -360 -7214
rect -1226 -7399 -1220 -7231
rect -1186 -7264 -1180 -7231
rect -316 -7231 -270 -7141
rect -316 -7264 -310 -7231
rect -1186 -7352 -310 -7264
rect -1186 -7399 -1180 -7352
rect -1226 -7411 -1180 -7399
rect -316 -7399 -310 -7352
rect -276 -7399 -270 -7231
rect -784 -7418 -684 -7408
rect -316 -7411 -270 -7399
rect -93 -7183 -41 -6509
rect -1148 -7427 -784 -7421
rect -684 -7427 -348 -7421
rect -1148 -7461 -1136 -7427
rect -360 -7461 -348 -7427
rect -1148 -7467 -784 -7461
rect -684 -7467 -348 -7461
rect -1226 -7489 -1180 -7477
rect -784 -7480 -684 -7470
rect -316 -7479 -270 -7477
rect -1226 -7657 -1220 -7489
rect -1186 -7529 -1180 -7489
rect -319 -7489 -267 -7479
rect -1186 -7549 -319 -7529
rect -1186 -7601 -783 -7549
rect -683 -7589 -319 -7549
rect -683 -7601 -310 -7589
rect -1186 -7617 -310 -7601
rect -1186 -7657 -1180 -7617
rect -1226 -7747 -1180 -7657
rect -316 -7657 -310 -7617
rect -276 -7599 -267 -7589
rect -276 -7657 -270 -7599
rect -1136 -7676 -936 -7666
rect -1148 -7725 -1136 -7679
rect -936 -7685 -348 -7679
rect -360 -7719 -348 -7685
rect -936 -7725 -348 -7719
rect -1136 -7738 -936 -7728
rect -1226 -7915 -1220 -7747
rect -1186 -7786 -1180 -7747
rect -316 -7747 -270 -7657
rect -316 -7786 -310 -7747
rect -1186 -7811 -310 -7786
rect -1186 -7863 -785 -7811
rect -685 -7863 -310 -7811
rect -1186 -7879 -310 -7863
rect -1186 -7915 -1180 -7879
rect -1226 -7927 -1180 -7915
rect -316 -7915 -310 -7879
rect -276 -7915 -270 -7747
rect -784 -7934 -684 -7924
rect -316 -7927 -270 -7915
rect -1148 -7943 -784 -7937
rect -684 -7943 -348 -7937
rect -1148 -7977 -1136 -7943
rect -360 -7977 -348 -7943
rect -1148 -7983 -784 -7977
rect -684 -7983 -348 -7977
rect -93 -7957 -41 -7283
rect -1226 -8005 -1180 -7993
rect -784 -7996 -684 -7986
rect -316 -7995 -270 -7993
rect -1226 -8173 -1220 -8005
rect -1186 -8044 -1180 -8005
rect -319 -8005 -267 -7995
rect -1186 -8131 -319 -8044
rect -267 -8131 -257 -8109
rect -1186 -8132 -310 -8131
rect -1186 -8173 -1180 -8132
rect -329 -8154 -310 -8132
rect -1226 -8263 -1180 -8173
rect -316 -8173 -310 -8154
rect -276 -8154 -257 -8131
rect -276 -8173 -270 -8154
rect -560 -8190 -360 -8180
rect -1148 -8201 -560 -8195
rect -1148 -8235 -1136 -8201
rect -1148 -8241 -560 -8235
rect -360 -8241 -348 -8195
rect -560 -8256 -360 -8246
rect -1226 -8431 -1220 -8263
rect -1186 -8303 -1180 -8263
rect -316 -8263 -270 -8173
rect -316 -8303 -310 -8263
rect -1186 -8391 -310 -8303
rect -1186 -8431 -1180 -8391
rect -1226 -8521 -1180 -8431
rect -316 -8431 -310 -8391
rect -276 -8431 -270 -8263
rect -1136 -8444 -936 -8434
rect -1148 -8499 -1136 -8453
rect -936 -8459 -348 -8453
rect -360 -8493 -348 -8459
rect -936 -8499 -348 -8493
rect -1136 -8518 -936 -8508
rect -1226 -8689 -1220 -8521
rect -1186 -8553 -1180 -8521
rect -316 -8521 -270 -8431
rect -316 -8553 -310 -8521
rect -1186 -8641 -310 -8553
rect -1186 -8689 -1180 -8641
rect -1226 -8779 -1180 -8689
rect -316 -8689 -310 -8641
rect -276 -8689 -270 -8521
rect -560 -8706 -360 -8696
rect -1148 -8717 -560 -8711
rect -1148 -8751 -1136 -8717
rect -1148 -8757 -560 -8751
rect -360 -8757 -348 -8711
rect -560 -8772 -360 -8762
rect -1226 -8947 -1220 -8779
rect -1186 -8816 -1180 -8779
rect -316 -8779 -270 -8689
rect -316 -8816 -310 -8779
rect -1186 -8904 -310 -8816
rect -1186 -8947 -1180 -8904
rect -1226 -8959 -1180 -8947
rect -316 -8947 -310 -8904
rect -276 -8947 -270 -8779
rect -784 -8966 -684 -8956
rect -316 -8959 -270 -8947
rect -93 -8731 -41 -8057
rect -1148 -8975 -784 -8969
rect -684 -8975 -348 -8969
rect -1148 -9009 -1136 -8975
rect -360 -9009 -348 -8975
rect -1148 -9015 -784 -9009
rect -684 -9015 -348 -9009
rect -1226 -9037 -1180 -9025
rect -784 -9028 -684 -9018
rect -316 -9027 -270 -9025
rect -1226 -9205 -1220 -9037
rect -1186 -9077 -1180 -9037
rect -319 -9037 -267 -9027
rect -1186 -9093 -319 -9077
rect -1186 -9145 -784 -9093
rect -684 -9137 -319 -9093
rect -684 -9145 -310 -9137
rect -1186 -9165 -310 -9145
rect -1186 -9205 -1180 -9165
rect -1226 -9295 -1180 -9205
rect -316 -9205 -310 -9165
rect -276 -9147 -267 -9137
rect -276 -9205 -270 -9147
rect -1136 -9224 -936 -9214
rect -1148 -9273 -1136 -9227
rect -936 -9233 -348 -9227
rect -360 -9267 -348 -9233
rect -936 -9273 -348 -9267
rect -1136 -9286 -936 -9276
rect -1226 -9463 -1220 -9295
rect -1186 -9340 -1180 -9295
rect -316 -9295 -270 -9205
rect -316 -9340 -310 -9295
rect -1186 -9358 -310 -9340
rect -1186 -9410 -784 -9358
rect -684 -9410 -310 -9358
rect -1186 -9429 -310 -9410
rect -1186 -9463 -1180 -9429
rect -1226 -9475 -1180 -9463
rect -316 -9463 -310 -9429
rect -276 -9463 -270 -9295
rect -784 -9482 -684 -9472
rect -316 -9475 -270 -9463
rect -1148 -9491 -784 -9485
rect -684 -9491 -348 -9485
rect -1148 -9525 -1136 -9491
rect -360 -9525 -348 -9491
rect -1148 -9531 -784 -9525
rect -684 -9531 -348 -9525
rect -93 -9505 -41 -8831
rect -1226 -9553 -1180 -9541
rect -784 -9544 -684 -9534
rect -316 -9543 -270 -9541
rect -1226 -9721 -1220 -9553
rect -1186 -9589 -1180 -9553
rect -319 -9553 -267 -9543
rect -1186 -9653 -319 -9589
rect -1186 -9678 -310 -9653
rect -1186 -9721 -1180 -9678
rect -1226 -9811 -1180 -9721
rect -316 -9721 -310 -9678
rect -276 -9663 -267 -9653
rect -276 -9721 -270 -9663
rect -560 -9738 -360 -9728
rect -1148 -9749 -560 -9743
rect -1148 -9783 -1136 -9749
rect -1148 -9789 -560 -9783
rect -360 -9789 -348 -9743
rect -560 -9804 -360 -9794
rect -1226 -9979 -1220 -9811
rect -1186 -9853 -1180 -9811
rect -316 -9811 -270 -9721
rect -316 -9853 -310 -9811
rect -1186 -9942 -310 -9853
rect -1186 -9979 -1180 -9942
rect -1226 -9991 -1180 -9979
rect -316 -9979 -310 -9942
rect -276 -9979 -270 -9811
rect -1136 -9992 -936 -9982
rect -316 -9991 -270 -9979
rect -1148 -10047 -1136 -10001
rect -936 -10007 -348 -10001
rect -360 -10041 -348 -10007
rect -936 -10047 -348 -10041
rect -1136 -10066 -936 -10056
rect -93 -10124 -41 -9605
rect 52 -3829 104 -3819
rect 333 -3849 345 -3815
rect 333 -3855 921 -3849
rect 1121 -3855 1133 -3809
rect 255 -3867 301 -3865
rect 52 -4345 104 -3929
rect 252 -3877 304 -3867
rect 921 -3868 1121 -3858
rect 1165 -3877 1211 -3865
rect 1165 -3918 1171 -3877
rect 304 -3938 1171 -3918
rect 304 -3977 644 -3938
rect 252 -3987 261 -3977
rect 255 -4045 261 -3987
rect 295 -3990 644 -3977
rect 744 -3990 1171 -3938
rect 295 -4006 1171 -3990
rect 295 -4045 301 -4006
rect 255 -4057 301 -4045
rect 1165 -4045 1171 -4006
rect 1205 -4045 1211 -3877
rect 646 -4064 746 -4054
rect 1165 -4057 1211 -4045
rect 333 -4073 646 -4067
rect 746 -4073 1133 -4067
rect 333 -4107 345 -4073
rect 1121 -4107 1133 -4073
rect 333 -4113 646 -4107
rect 746 -4113 1133 -4107
rect 255 -4125 301 -4123
rect 252 -4135 304 -4125
rect 646 -4126 746 -4116
rect 1165 -4135 1211 -4123
rect 1165 -4171 1171 -4135
rect 304 -4259 1171 -4171
rect 1165 -4303 1171 -4259
rect 1205 -4303 1211 -4135
rect 252 -4329 304 -4319
rect 921 -4320 1121 -4310
rect 52 -5119 104 -4445
rect 255 -4393 301 -4329
rect 333 -4331 921 -4325
rect 333 -4365 345 -4331
rect 333 -4371 921 -4365
rect 1121 -4371 1133 -4325
rect 921 -4386 1121 -4376
rect 255 -4561 261 -4393
rect 295 -4431 301 -4393
rect 1165 -4393 1211 -4303
rect 1165 -4431 1171 -4393
rect 295 -4519 1171 -4431
rect 295 -4561 301 -4519
rect 255 -4651 301 -4561
rect 1165 -4561 1171 -4519
rect 1205 -4561 1211 -4393
rect 345 -4574 545 -4564
rect 333 -4629 345 -4583
rect 545 -4589 1133 -4583
rect 1121 -4623 1133 -4589
rect 545 -4629 1133 -4623
rect 345 -4648 545 -4638
rect 255 -4819 261 -4651
rect 295 -4690 301 -4651
rect 1165 -4651 1211 -4561
rect 1165 -4690 1171 -4651
rect 295 -4778 1171 -4690
rect 295 -4819 301 -4778
rect 255 -4909 301 -4819
rect 1165 -4819 1171 -4778
rect 1205 -4819 1211 -4651
rect 921 -4836 1121 -4826
rect 333 -4847 921 -4841
rect 333 -4881 345 -4847
rect 333 -4887 921 -4881
rect 1121 -4887 1133 -4841
rect 921 -4902 1121 -4892
rect 255 -5077 261 -4909
rect 295 -4946 301 -4909
rect 1165 -4909 1211 -4819
rect 1165 -4946 1171 -4909
rect 295 -5034 1171 -4946
rect 295 -5077 301 -5034
rect 255 -5089 301 -5077
rect 1165 -5077 1171 -5034
rect 1205 -5077 1211 -4909
rect 646 -5096 746 -5086
rect 1165 -5089 1211 -5077
rect 333 -5105 646 -5099
rect 746 -5105 1133 -5099
rect 333 -5139 345 -5105
rect 1121 -5139 1133 -5105
rect 333 -5145 646 -5139
rect 746 -5145 1133 -5139
rect 255 -5157 301 -5155
rect 52 -5893 104 -5219
rect 252 -5167 304 -5157
rect 646 -5158 746 -5148
rect 1165 -5167 1211 -5155
rect 1165 -5198 1171 -5167
rect 304 -5230 1171 -5198
rect 304 -5267 646 -5230
rect 252 -5277 261 -5267
rect 255 -5335 261 -5277
rect 295 -5282 646 -5267
rect 746 -5282 1171 -5230
rect 295 -5304 1171 -5282
rect 295 -5335 301 -5304
rect 255 -5425 301 -5335
rect 1165 -5335 1171 -5304
rect 1205 -5335 1211 -5167
rect 921 -5354 1121 -5344
rect 333 -5363 921 -5357
rect 333 -5397 345 -5363
rect 333 -5403 921 -5397
rect 1121 -5403 1133 -5357
rect 921 -5416 1121 -5406
rect 255 -5593 261 -5425
rect 295 -5453 301 -5425
rect 1165 -5425 1211 -5335
rect 1165 -5453 1171 -5425
rect 295 -5485 1171 -5453
rect 295 -5537 648 -5485
rect 748 -5537 1171 -5485
rect 295 -5559 1171 -5537
rect 295 -5593 301 -5559
rect 255 -5605 301 -5593
rect 1165 -5593 1171 -5559
rect 1205 -5593 1211 -5425
rect 646 -5612 746 -5602
rect 1165 -5605 1211 -5593
rect 333 -5621 646 -5615
rect 746 -5621 1133 -5615
rect 333 -5655 345 -5621
rect 1121 -5655 1133 -5621
rect 333 -5661 646 -5655
rect 746 -5661 1133 -5655
rect 255 -5673 301 -5671
rect 252 -5683 304 -5673
rect 646 -5674 746 -5664
rect 1165 -5683 1211 -5671
rect 1165 -5726 1171 -5683
rect 304 -5814 1171 -5726
rect 1165 -5851 1171 -5814
rect 1205 -5851 1211 -5683
rect 252 -5877 304 -5867
rect 921 -5868 1121 -5858
rect 52 -6667 104 -5993
rect 255 -5941 301 -5877
rect 333 -5879 921 -5873
rect 333 -5913 345 -5879
rect 333 -5919 921 -5913
rect 1121 -5919 1133 -5873
rect 921 -5934 1121 -5924
rect 255 -6109 261 -5941
rect 295 -5981 301 -5941
rect 1165 -5941 1211 -5851
rect 1165 -5981 1171 -5941
rect 295 -6069 1171 -5981
rect 295 -6109 301 -6069
rect 255 -6199 301 -6109
rect 1165 -6109 1171 -6069
rect 1205 -6109 1211 -5941
rect 345 -6122 545 -6112
rect 333 -6177 345 -6131
rect 545 -6137 1133 -6131
rect 1121 -6171 1133 -6137
rect 545 -6177 1133 -6171
rect 345 -6196 545 -6186
rect 255 -6367 261 -6199
rect 295 -6242 301 -6199
rect 1165 -6199 1211 -6109
rect 1165 -6242 1171 -6199
rect 295 -6330 1171 -6242
rect 295 -6367 301 -6330
rect 255 -6457 301 -6367
rect 1165 -6367 1171 -6330
rect 1205 -6367 1211 -6199
rect 921 -6384 1121 -6374
rect 333 -6395 921 -6389
rect 333 -6429 345 -6395
rect 333 -6435 921 -6429
rect 1121 -6435 1133 -6389
rect 921 -6450 1121 -6440
rect 255 -6625 261 -6457
rect 295 -6498 301 -6457
rect 1165 -6457 1211 -6367
rect 1165 -6498 1171 -6457
rect 295 -6586 1171 -6498
rect 295 -6625 301 -6586
rect 255 -6637 301 -6625
rect 1165 -6625 1171 -6586
rect 1205 -6625 1211 -6457
rect 645 -6644 745 -6634
rect 1165 -6637 1211 -6625
rect 333 -6653 645 -6647
rect 745 -6653 1133 -6647
rect 333 -6687 345 -6653
rect 1121 -6687 1133 -6653
rect 333 -6693 645 -6687
rect 745 -6693 1133 -6687
rect 255 -6705 301 -6703
rect 52 -7441 104 -6767
rect 252 -6715 304 -6705
rect 645 -6706 745 -6696
rect 1165 -6715 1211 -6703
rect 1165 -6767 1171 -6715
rect 304 -6781 1171 -6767
rect 304 -6815 648 -6781
rect 252 -6825 261 -6815
rect 255 -6883 261 -6825
rect 295 -6833 648 -6815
rect 748 -6833 1171 -6781
rect 295 -6848 1171 -6833
rect 295 -6883 301 -6848
rect 255 -6973 301 -6883
rect 1165 -6883 1171 -6848
rect 1205 -6883 1211 -6715
rect 921 -6902 1121 -6892
rect 333 -6911 921 -6905
rect 333 -6945 345 -6911
rect 333 -6951 921 -6945
rect 1121 -6951 1133 -6905
rect 921 -6964 1121 -6954
rect 255 -7141 261 -6973
rect 295 -7027 301 -6973
rect 1165 -6973 1211 -6883
rect 1165 -7027 1171 -6973
rect 295 -7043 1171 -7027
rect 295 -7095 646 -7043
rect 746 -7095 1171 -7043
rect 295 -7108 1171 -7095
rect 295 -7141 301 -7108
rect 255 -7153 301 -7141
rect 1165 -7141 1171 -7108
rect 1205 -7141 1211 -6973
rect 646 -7160 746 -7150
rect 1165 -7153 1211 -7141
rect 333 -7169 646 -7163
rect 746 -7169 1133 -7163
rect 333 -7203 345 -7169
rect 1121 -7203 1133 -7169
rect 333 -7209 646 -7203
rect 746 -7209 1133 -7203
rect 255 -7221 301 -7219
rect 252 -7231 304 -7221
rect 646 -7222 746 -7212
rect 1165 -7231 1211 -7219
rect 1165 -7266 1171 -7231
rect 304 -7354 1171 -7266
rect 1165 -7399 1171 -7354
rect 1205 -7399 1211 -7231
rect 252 -7425 304 -7415
rect 921 -7416 1121 -7406
rect 52 -8215 104 -7541
rect 255 -7489 301 -7425
rect 333 -7427 921 -7421
rect 333 -7461 345 -7427
rect 333 -7467 921 -7461
rect 1121 -7467 1133 -7421
rect 921 -7482 1121 -7472
rect 255 -7657 261 -7489
rect 295 -7537 301 -7489
rect 1165 -7489 1211 -7399
rect 1165 -7537 1171 -7489
rect 295 -7625 1171 -7537
rect 295 -7657 301 -7625
rect 255 -7747 301 -7657
rect 1165 -7657 1171 -7625
rect 1205 -7657 1211 -7489
rect 345 -7670 545 -7660
rect 333 -7725 345 -7679
rect 545 -7685 1133 -7679
rect 1121 -7719 1133 -7685
rect 545 -7725 1133 -7719
rect 345 -7744 545 -7734
rect 255 -7915 261 -7747
rect 295 -7789 301 -7747
rect 1165 -7747 1211 -7657
rect 1165 -7789 1171 -7747
rect 295 -7877 1171 -7789
rect 295 -7915 301 -7877
rect 255 -8005 301 -7915
rect 1165 -7915 1171 -7877
rect 1205 -7915 1211 -7747
rect 921 -7932 1121 -7922
rect 333 -7943 921 -7937
rect 333 -7977 345 -7943
rect 333 -7983 921 -7977
rect 1121 -7983 1133 -7937
rect 921 -7998 1121 -7988
rect 255 -8173 261 -8005
rect 295 -8042 301 -8005
rect 1165 -8005 1211 -7915
rect 1165 -8042 1171 -8005
rect 295 -8130 1171 -8042
rect 295 -8173 301 -8130
rect 255 -8185 301 -8173
rect 1165 -8173 1171 -8130
rect 1205 -8173 1211 -8005
rect 646 -8192 746 -8182
rect 1165 -8185 1211 -8173
rect 333 -8201 646 -8195
rect 746 -8201 1133 -8195
rect 333 -8235 345 -8201
rect 1121 -8235 1133 -8201
rect 333 -8241 646 -8235
rect 746 -8241 1133 -8235
rect 255 -8253 301 -8251
rect 52 -8989 104 -8315
rect 252 -8263 304 -8253
rect 646 -8254 746 -8244
rect 1165 -8263 1211 -8251
rect 1165 -8309 1171 -8263
rect 304 -8329 1171 -8309
rect 304 -8363 644 -8329
rect 252 -8373 261 -8363
rect 255 -8431 261 -8373
rect 295 -8381 644 -8363
rect 744 -8381 1171 -8329
rect 295 -8397 1171 -8381
rect 295 -8431 301 -8397
rect 255 -8521 301 -8431
rect 1165 -8431 1171 -8397
rect 1205 -8431 1211 -8263
rect 921 -8450 1121 -8440
rect 333 -8459 921 -8453
rect 333 -8493 345 -8459
rect 333 -8499 921 -8493
rect 1121 -8499 1133 -8453
rect 921 -8512 1121 -8502
rect 255 -8689 261 -8521
rect 295 -8563 301 -8521
rect 1165 -8521 1211 -8431
rect 1165 -8563 1171 -8521
rect 295 -8585 1171 -8563
rect 295 -8637 645 -8585
rect 745 -8637 1171 -8585
rect 295 -8651 1171 -8637
rect 295 -8689 301 -8651
rect 255 -8701 301 -8689
rect 1165 -8689 1171 -8651
rect 1205 -8689 1211 -8521
rect 646 -8708 746 -8698
rect 1165 -8701 1211 -8689
rect 333 -8717 646 -8711
rect 746 -8717 1133 -8711
rect 333 -8751 345 -8717
rect 1121 -8751 1133 -8717
rect 333 -8757 646 -8751
rect 746 -8757 1133 -8751
rect 255 -8769 301 -8767
rect 252 -8779 304 -8769
rect 646 -8770 746 -8760
rect 1165 -8779 1211 -8767
rect 1165 -8826 1171 -8779
rect 304 -8914 1171 -8826
rect 1165 -8947 1171 -8914
rect 1205 -8947 1211 -8779
rect 921 -8964 1121 -8954
rect 252 -8989 304 -8979
rect 333 -8975 921 -8969
rect 52 -9763 104 -9089
rect 255 -9037 301 -8989
rect 333 -9009 345 -8975
rect 333 -9015 921 -9009
rect 1121 -9015 1133 -8969
rect 921 -9030 1121 -9020
rect 255 -9205 261 -9037
rect 295 -9075 301 -9037
rect 1165 -9037 1211 -8947
rect 1165 -9075 1171 -9037
rect 295 -9163 1171 -9075
rect 295 -9205 301 -9163
rect 255 -9295 301 -9205
rect 1165 -9205 1171 -9163
rect 1205 -9205 1211 -9037
rect 345 -9218 545 -9208
rect 333 -9273 345 -9227
rect 545 -9233 1133 -9227
rect 1121 -9267 1133 -9233
rect 545 -9273 1133 -9267
rect 345 -9292 545 -9282
rect 255 -9463 261 -9295
rect 295 -9345 301 -9295
rect 1165 -9295 1211 -9205
rect 1165 -9345 1171 -9295
rect 295 -9433 1171 -9345
rect 295 -9463 301 -9433
rect 255 -9553 301 -9463
rect 1165 -9463 1171 -9433
rect 1205 -9463 1211 -9295
rect 920 -9480 1120 -9470
rect 333 -9491 920 -9485
rect 1120 -9491 1133 -9485
rect 333 -9525 345 -9491
rect 1121 -9525 1133 -9491
rect 333 -9531 920 -9525
rect 1120 -9531 1133 -9525
rect 920 -9546 1120 -9536
rect 255 -9721 261 -9553
rect 295 -9594 301 -9553
rect 1165 -9553 1211 -9463
rect 1165 -9594 1171 -9553
rect 295 -9682 1171 -9594
rect 295 -9721 301 -9682
rect 255 -9733 301 -9721
rect 1165 -9721 1171 -9682
rect 1205 -9721 1211 -9553
rect 646 -9740 746 -9730
rect 1165 -9733 1211 -9721
rect 333 -9749 646 -9743
rect 746 -9749 1133 -9743
rect 333 -9783 345 -9749
rect 1121 -9783 1133 -9749
rect 333 -9789 646 -9783
rect 746 -9789 1133 -9783
rect 255 -9801 301 -9799
rect 52 -9985 104 -9863
rect 252 -9811 304 -9801
rect 646 -9802 746 -9792
rect 1165 -9811 1211 -9799
rect 1165 -9846 1171 -9811
rect 304 -9863 1171 -9846
rect 304 -9911 648 -9863
rect 252 -9921 261 -9911
rect 255 -9979 261 -9921
rect 295 -9915 648 -9911
rect 748 -9915 1171 -9863
rect 295 -9934 1171 -9915
rect 295 -9979 301 -9934
rect 255 -9991 301 -9979
rect 1165 -9979 1171 -9934
rect 1205 -9979 1211 -9811
rect 921 -9998 1121 -9988
rect 1165 -9991 1211 -9979
rect 333 -10007 921 -10001
rect 333 -10041 345 -10007
rect 333 -10047 921 -10041
rect 1121 -10047 1133 -10001
rect 921 -10060 1121 -10050
rect 1374 -10070 1380 -3729
rect 1492 -10070 1498 -3729
rect 2116 -8325 2122 -2918
rect 2313 -8325 2319 -2918
rect 3269 -2936 3392 -2926
rect 3257 -2985 3269 -2939
rect 3392 -2945 3457 -2939
rect 3445 -2979 3457 -2945
rect 3392 -2985 3457 -2979
rect 2482 -3001 2542 -2991
rect 2470 -3050 2482 -3004
rect 2598 -3001 2658 -2991
rect 2542 -3010 2598 -3004
rect 2542 -3050 2598 -3044
rect 2392 -3072 2438 -3060
rect 2482 -3063 2542 -3053
rect 2658 -3050 2670 -3004
rect 3170 -3007 3216 -2990
rect 3269 -2998 3392 -2988
rect 2598 -3063 2658 -3053
rect 2392 -3240 2398 -3072
rect 2432 -3114 2438 -3072
rect 2702 -3072 2748 -3060
rect 2702 -3114 2708 -3072
rect 2432 -3181 2708 -3114
rect 2432 -3240 2438 -3181
rect 2392 -3262 2438 -3240
rect 2702 -3240 2708 -3181
rect 2742 -3240 2748 -3072
rect 2702 -3249 2748 -3240
rect 2598 -3259 2748 -3249
rect 2392 -3268 2598 -3262
rect 2392 -3302 2482 -3268
rect 2392 -3308 2598 -3302
rect 2392 -3330 2438 -3308
rect 2658 -3311 2748 -3259
rect 2598 -3321 2748 -3311
rect 2392 -3498 2398 -3330
rect 2432 -3381 2438 -3330
rect 2702 -3330 2748 -3321
rect 2702 -3381 2708 -3330
rect 2432 -3448 2708 -3381
rect 2432 -3498 2438 -3448
rect 2392 -3588 2438 -3498
rect 2702 -3498 2708 -3448
rect 2742 -3498 2748 -3330
rect 2482 -3517 2542 -3507
rect 2470 -3566 2482 -3520
rect 2542 -3526 2670 -3520
rect 2658 -3560 2670 -3526
rect 2542 -3566 2670 -3560
rect 2482 -3579 2542 -3569
rect 2392 -3756 2398 -3588
rect 2432 -3640 2438 -3588
rect 2702 -3588 2748 -3498
rect 2702 -3640 2708 -3588
rect 2432 -3707 2708 -3640
rect 2432 -3756 2438 -3707
rect 2392 -3778 2438 -3756
rect 2702 -3756 2708 -3707
rect 2742 -3756 2748 -3588
rect 2702 -3765 2748 -3756
rect 2598 -3775 2748 -3765
rect 2392 -3784 2598 -3778
rect 2392 -3818 2482 -3784
rect 2392 -3824 2598 -3818
rect 2392 -3846 2438 -3824
rect 2658 -3827 2748 -3775
rect 2598 -3837 2748 -3827
rect 2392 -4014 2398 -3846
rect 2432 -3900 2438 -3846
rect 2702 -3846 2748 -3837
rect 2702 -3900 2708 -3846
rect 2432 -3967 2708 -3900
rect 2432 -4014 2438 -3967
rect 2392 -4104 2438 -4014
rect 2702 -4014 2708 -3967
rect 2742 -4014 2748 -3846
rect 2482 -4033 2542 -4023
rect 2470 -4082 2482 -4036
rect 2542 -4042 2670 -4036
rect 2658 -4076 2670 -4042
rect 2542 -4082 2670 -4076
rect 2482 -4095 2542 -4085
rect 2392 -4272 2398 -4104
rect 2432 -4162 2438 -4104
rect 2702 -4104 2748 -4014
rect 2702 -4162 2708 -4104
rect 2432 -4229 2708 -4162
rect 2432 -4272 2438 -4229
rect 2392 -4284 2438 -4272
rect 2702 -4272 2708 -4229
rect 2742 -4272 2748 -4104
rect 2482 -4291 2542 -4281
rect 2702 -4284 2748 -4272
rect 3170 -3375 3176 -3007
rect 3210 -3044 3216 -3007
rect 3498 -3007 3544 -2995
rect 3498 -3044 3504 -3007
rect 3210 -3323 3504 -3044
rect 3210 -3375 3216 -3323
rect 3170 -3588 3216 -3375
rect 3498 -3375 3504 -3323
rect 3538 -3375 3544 -3007
rect 3322 -3394 3445 -3384
rect 3498 -3387 3544 -3375
rect 3257 -3403 3322 -3397
rect 3257 -3437 3269 -3403
rect 3257 -3443 3322 -3437
rect 3445 -3443 3457 -3397
rect 3322 -3456 3445 -3446
rect 3269 -3517 3392 -3507
rect 3257 -3566 3269 -3520
rect 3392 -3526 3457 -3520
rect 3445 -3560 3457 -3526
rect 3392 -3566 3457 -3560
rect 3269 -3579 3392 -3569
rect 3170 -3956 3176 -3588
rect 3210 -3620 3216 -3588
rect 3498 -3588 3544 -3576
rect 3498 -3620 3504 -3588
rect 3210 -3899 3504 -3620
rect 3210 -3956 3216 -3899
rect 2470 -4340 2482 -4294
rect 2542 -4300 2670 -4294
rect 2658 -4334 2670 -4300
rect 2542 -4340 2670 -4334
rect 2392 -4362 2438 -4350
rect 2482 -4353 2542 -4343
rect 2392 -4530 2398 -4362
rect 2432 -4422 2438 -4362
rect 2702 -4362 2748 -4350
rect 2702 -4422 2708 -4362
rect 2432 -4489 2708 -4422
rect 2432 -4530 2438 -4489
rect 2392 -4552 2438 -4530
rect 2702 -4530 2708 -4489
rect 2742 -4530 2748 -4362
rect 2702 -4539 2748 -4530
rect 2598 -4549 2748 -4539
rect 2392 -4558 2598 -4552
rect 2392 -4592 2482 -4558
rect 2392 -4598 2598 -4592
rect 2392 -4620 2438 -4598
rect 2658 -4601 2748 -4549
rect 2598 -4611 2748 -4601
rect 2392 -4788 2398 -4620
rect 2432 -4672 2438 -4620
rect 2702 -4620 2748 -4611
rect 2702 -4672 2708 -4620
rect 2432 -4739 2708 -4672
rect 2432 -4788 2438 -4739
rect 2392 -4878 2438 -4788
rect 2702 -4788 2708 -4739
rect 2742 -4788 2748 -4620
rect 2482 -4807 2542 -4797
rect 2470 -4856 2482 -4810
rect 2542 -4816 2670 -4810
rect 2658 -4850 2670 -4816
rect 2542 -4856 2670 -4850
rect 2482 -4869 2542 -4859
rect 2392 -5046 2398 -4878
rect 2432 -4931 2438 -4878
rect 2702 -4878 2748 -4788
rect 2702 -4931 2708 -4878
rect 2432 -4998 2708 -4931
rect 2432 -5046 2438 -4998
rect 2392 -5068 2438 -5046
rect 2702 -5046 2708 -4998
rect 2742 -5046 2748 -4878
rect 2702 -5055 2748 -5046
rect 2598 -5065 2748 -5055
rect 2392 -5074 2598 -5068
rect 2392 -5108 2482 -5074
rect 2392 -5114 2598 -5108
rect 2392 -5136 2438 -5114
rect 2658 -5117 2748 -5065
rect 2598 -5127 2748 -5117
rect 2392 -5304 2398 -5136
rect 2432 -5192 2438 -5136
rect 2702 -5136 2748 -5127
rect 2702 -5192 2708 -5136
rect 2432 -5259 2708 -5192
rect 2432 -5304 2438 -5259
rect 2392 -5394 2438 -5304
rect 2702 -5304 2708 -5259
rect 2742 -5304 2748 -5136
rect 2482 -5323 2542 -5313
rect 2470 -5372 2482 -5326
rect 2542 -5332 2670 -5326
rect 2658 -5366 2670 -5332
rect 2542 -5372 2670 -5366
rect 2482 -5385 2542 -5375
rect 2392 -5562 2398 -5394
rect 2432 -5449 2438 -5394
rect 2702 -5394 2748 -5304
rect 2702 -5449 2708 -5394
rect 2432 -5516 2708 -5449
rect 2432 -5562 2438 -5516
rect 2392 -5574 2438 -5562
rect 2702 -5562 2708 -5516
rect 2742 -5562 2748 -5394
rect 2482 -5581 2542 -5571
rect 2702 -5574 2748 -5562
rect 3170 -4878 3216 -3956
rect 3498 -3956 3504 -3899
rect 3538 -3956 3544 -3588
rect 3321 -3975 3445 -3965
rect 3498 -3968 3544 -3956
rect 3257 -3984 3321 -3978
rect 3257 -4018 3269 -3984
rect 3257 -4024 3321 -4018
rect 3445 -4024 3457 -3978
rect 3321 -4037 3445 -4027
rect 3706 -4215 3710 -4157
rect 3269 -4807 3382 -4797
rect 3257 -4856 3269 -4810
rect 3382 -4816 3457 -4810
rect 3445 -4850 3457 -4816
rect 3382 -4856 3457 -4850
rect 3269 -4869 3382 -4859
rect 3170 -5246 3176 -4878
rect 3210 -4930 3216 -4878
rect 3498 -4878 3544 -4866
rect 3498 -4930 3504 -4878
rect 3210 -5209 3504 -4930
rect 3210 -5246 3216 -5209
rect 2470 -5630 2482 -5584
rect 2542 -5590 2670 -5584
rect 2658 -5624 2670 -5590
rect 2542 -5630 2670 -5624
rect 2392 -5652 2438 -5640
rect 2482 -5643 2542 -5633
rect 2392 -5820 2398 -5652
rect 2432 -5707 2438 -5652
rect 2702 -5652 2748 -5640
rect 2702 -5707 2708 -5652
rect 2432 -5774 2708 -5707
rect 2432 -5820 2438 -5774
rect 2392 -5842 2438 -5820
rect 2702 -5820 2708 -5774
rect 2742 -5820 2748 -5652
rect 2702 -5829 2748 -5820
rect 2598 -5839 2748 -5829
rect 2392 -5848 2598 -5842
rect 2392 -5882 2482 -5848
rect 2392 -5888 2598 -5882
rect 2392 -5910 2438 -5888
rect 2658 -5891 2748 -5839
rect 2598 -5901 2748 -5891
rect 2392 -6078 2398 -5910
rect 2432 -5969 2438 -5910
rect 2702 -5910 2748 -5901
rect 2702 -5969 2708 -5910
rect 2432 -6036 2708 -5969
rect 2432 -6078 2438 -6036
rect 2392 -6168 2438 -6078
rect 2702 -6078 2708 -6036
rect 2742 -6078 2748 -5910
rect 2482 -6097 2542 -6087
rect 2470 -6146 2482 -6100
rect 2542 -6106 2670 -6100
rect 2658 -6140 2670 -6106
rect 2542 -6146 2670 -6140
rect 2482 -6159 2542 -6149
rect 2392 -6336 2398 -6168
rect 2432 -6222 2438 -6168
rect 2702 -6168 2748 -6078
rect 2702 -6222 2708 -6168
rect 2432 -6289 2708 -6222
rect 2432 -6336 2438 -6289
rect 2392 -6358 2438 -6336
rect 2702 -6336 2708 -6289
rect 2742 -6336 2748 -6168
rect 2702 -6345 2748 -6336
rect 2598 -6355 2748 -6345
rect 2392 -6364 2598 -6358
rect 2392 -6398 2482 -6364
rect 2392 -6404 2598 -6398
rect 2392 -6426 2438 -6404
rect 2658 -6407 2748 -6355
rect 2598 -6417 2748 -6407
rect 2392 -6594 2398 -6426
rect 2432 -6483 2438 -6426
rect 2702 -6426 2748 -6417
rect 2702 -6483 2708 -6426
rect 2432 -6550 2708 -6483
rect 2432 -6594 2438 -6550
rect 2392 -6684 2438 -6594
rect 2702 -6594 2708 -6550
rect 2742 -6594 2748 -6426
rect 2482 -6613 2542 -6603
rect 2470 -6662 2482 -6616
rect 2542 -6622 2670 -6616
rect 2658 -6656 2670 -6622
rect 2542 -6662 2670 -6656
rect 2482 -6675 2542 -6665
rect 2392 -6852 2398 -6684
rect 2432 -6737 2438 -6684
rect 2702 -6684 2748 -6594
rect 2702 -6737 2708 -6684
rect 2432 -6804 2708 -6737
rect 2432 -6852 2438 -6804
rect 2392 -6864 2438 -6852
rect 2702 -6852 2708 -6804
rect 2742 -6852 2748 -6684
rect 2482 -6871 2542 -6861
rect 2702 -6864 2748 -6852
rect 3170 -6168 3216 -5246
rect 3498 -5246 3504 -5209
rect 3538 -5246 3544 -4878
rect 3322 -5265 3445 -5255
rect 3498 -5258 3544 -5246
rect 3257 -5274 3322 -5268
rect 3257 -5308 3269 -5274
rect 3257 -5314 3322 -5308
rect 3445 -5314 3457 -5268
rect 3322 -5327 3445 -5317
rect 3269 -6097 3382 -6087
rect 3257 -6146 3269 -6100
rect 3382 -6106 3457 -6100
rect 3445 -6140 3457 -6106
rect 3382 -6146 3457 -6140
rect 3269 -6159 3382 -6149
rect 3170 -6536 3176 -6168
rect 3210 -6211 3216 -6168
rect 3498 -6168 3544 -6156
rect 3498 -6211 3504 -6168
rect 3210 -6490 3504 -6211
rect 3210 -6536 3216 -6490
rect 2470 -6920 2482 -6874
rect 2542 -6880 2670 -6874
rect 2658 -6914 2670 -6880
rect 2542 -6920 2670 -6914
rect 2392 -6942 2438 -6930
rect 2482 -6933 2542 -6923
rect 2392 -7110 2398 -6942
rect 2432 -6989 2438 -6942
rect 2702 -6942 2748 -6930
rect 2702 -6989 2708 -6942
rect 2432 -7056 2708 -6989
rect 2432 -7110 2438 -7056
rect 2392 -7132 2438 -7110
rect 2702 -7110 2708 -7056
rect 2742 -7110 2748 -6942
rect 2702 -7119 2748 -7110
rect 2598 -7129 2748 -7119
rect 2392 -7138 2598 -7132
rect 2392 -7172 2482 -7138
rect 2392 -7178 2598 -7172
rect 2392 -7200 2438 -7178
rect 2658 -7181 2748 -7129
rect 2598 -7191 2748 -7181
rect 2392 -7368 2398 -7200
rect 2432 -7249 2438 -7200
rect 2702 -7200 2748 -7191
rect 2702 -7249 2708 -7200
rect 2432 -7316 2708 -7249
rect 2432 -7368 2438 -7316
rect 2392 -7458 2438 -7368
rect 2702 -7368 2708 -7316
rect 2742 -7368 2748 -7200
rect 2482 -7387 2542 -7377
rect 2470 -7436 2482 -7390
rect 2542 -7396 2670 -7390
rect 2658 -7430 2670 -7396
rect 2542 -7436 2670 -7430
rect 2482 -7449 2542 -7439
rect 2392 -7626 2398 -7458
rect 2432 -7506 2438 -7458
rect 2702 -7458 2748 -7368
rect 2702 -7506 2708 -7458
rect 2432 -7573 2708 -7506
rect 2432 -7626 2438 -7573
rect 2392 -7648 2438 -7626
rect 2702 -7626 2708 -7573
rect 2742 -7626 2748 -7458
rect 2702 -7635 2748 -7626
rect 2598 -7645 2748 -7635
rect 2392 -7654 2598 -7648
rect 2392 -7688 2482 -7654
rect 2392 -7694 2598 -7688
rect 2392 -7716 2438 -7694
rect 2658 -7697 2748 -7645
rect 2598 -7707 2748 -7697
rect 2392 -7884 2398 -7716
rect 2432 -7768 2438 -7716
rect 2702 -7716 2748 -7707
rect 2702 -7768 2708 -7716
rect 2432 -7835 2708 -7768
rect 2432 -7884 2438 -7835
rect 2392 -7974 2438 -7884
rect 2702 -7884 2708 -7835
rect 2742 -7884 2748 -7716
rect 2482 -7903 2542 -7893
rect 2470 -7952 2482 -7906
rect 2542 -7912 2670 -7906
rect 2658 -7946 2670 -7912
rect 2542 -7952 2670 -7946
rect 2482 -7965 2542 -7955
rect 2392 -8142 2398 -7974
rect 2432 -8026 2438 -7974
rect 2702 -7974 2748 -7884
rect 2702 -8026 2708 -7974
rect 2432 -8093 2708 -8026
rect 2432 -8142 2438 -8093
rect 2392 -8154 2438 -8142
rect 2702 -8142 2708 -8093
rect 2742 -8142 2748 -7974
rect 2482 -8161 2542 -8151
rect 2702 -8154 2748 -8142
rect 3170 -7458 3216 -6536
rect 3498 -6536 3504 -6490
rect 3538 -6536 3544 -6168
rect 3322 -6555 3445 -6545
rect 3498 -6548 3544 -6536
rect 3257 -6564 3322 -6558
rect 3257 -6598 3269 -6564
rect 3257 -6604 3322 -6598
rect 3445 -6604 3457 -6558
rect 3322 -6617 3445 -6607
rect 3269 -7387 3382 -7377
rect 3257 -7436 3269 -7390
rect 3382 -7396 3457 -7390
rect 3445 -7430 3457 -7396
rect 3382 -7436 3457 -7430
rect 3269 -7449 3382 -7439
rect 3170 -7826 3176 -7458
rect 3210 -7509 3216 -7458
rect 3498 -7458 3544 -7446
rect 3498 -7509 3504 -7458
rect 3210 -7788 3504 -7509
rect 3210 -7826 3216 -7788
rect 2470 -8210 2482 -8164
rect 2542 -8170 2670 -8164
rect 2658 -8204 2670 -8170
rect 2542 -8210 2670 -8204
rect 2482 -8223 2542 -8213
rect 2116 -8337 2319 -8325
rect 3170 -8546 3216 -7826
rect 3498 -7826 3504 -7788
rect 3538 -7826 3544 -7458
rect 3322 -7845 3445 -7835
rect 3498 -7838 3544 -7826
rect 3257 -7854 3322 -7848
rect 3257 -7888 3269 -7854
rect 3257 -7894 3322 -7888
rect 3445 -7894 3457 -7848
rect 3322 -7907 3445 -7897
rect 3710 -7895 3716 -4242
rect 8442 -3760 8452 -2333
rect 9795 -2509 10341 -2503
rect 9795 -2510 9805 -2509
rect 8790 -3513 8800 -2510
rect 9709 -2629 9719 -2619
rect 9040 -2635 9719 -2629
rect 10128 -2629 10138 -2619
rect 9040 -2669 9052 -2635
rect 9040 -2675 9719 -2669
rect 9709 -2684 9719 -2675
rect 10128 -2675 10140 -2629
rect 10128 -2684 10138 -2675
rect 8962 -2697 9008 -2685
rect 8962 -2712 8968 -2697
rect 9002 -2712 9008 -2697
rect 10172 -2697 10218 -2685
rect 8947 -2852 8957 -2712
rect 9013 -2852 9023 -2712
rect 8962 -2965 8968 -2852
rect 9002 -2965 9008 -2852
rect 8962 -3055 9008 -2965
rect 10172 -2965 10178 -2697
rect 10212 -2965 10218 -2697
rect 9042 -2987 9052 -2978
rect 9040 -3033 9052 -2987
rect 9552 -2987 9562 -2978
rect 9552 -2993 10140 -2987
rect 10128 -3027 10140 -2993
rect 9042 -3042 9052 -3033
rect 9552 -3033 10140 -3027
rect 9552 -3042 9562 -3033
rect 8962 -3323 8968 -3055
rect 9002 -3323 9008 -3055
rect 8962 -3335 9008 -3323
rect 10172 -3055 10218 -2965
rect 10172 -3323 10178 -3055
rect 10212 -3323 10218 -3055
rect 10172 -3335 10218 -3323
rect 9709 -3345 9719 -3335
rect 9040 -3351 9719 -3345
rect 10128 -3345 10138 -3335
rect 9040 -3385 9052 -3351
rect 9040 -3391 9719 -3385
rect 9709 -3400 9719 -3391
rect 10128 -3391 10140 -3345
rect 10128 -3400 10138 -3391
rect 10331 -3513 10341 -2509
rect 8790 -3519 10341 -3513
rect 11117 -2503 11123 -2163
rect 11283 -2379 11293 -2377
rect 11281 -2429 11293 -2379
rect 11495 -2379 11505 -2377
rect 12117 -2379 12127 -2378
rect 11495 -2385 11702 -2379
rect 11690 -2423 11702 -2385
rect 11495 -2429 11702 -2423
rect 11920 -2385 12127 -2379
rect 12329 -2379 12339 -2378
rect 11920 -2423 11932 -2385
rect 11920 -2429 12127 -2423
rect 12117 -2430 12127 -2429
rect 12329 -2429 12341 -2379
rect 12329 -2430 12339 -2429
rect 10552 -2509 11123 -2503
rect 8679 -3760 10341 -3758
rect 8446 -3764 10341 -3760
rect 8446 -3772 8685 -3764
rect 10331 -3769 10341 -3764
rect 10552 -3769 10562 -2509
rect 10922 -2515 11123 -2509
rect 10335 -3781 10558 -3769
rect 3861 -4215 3865 -4157
rect 3855 -7895 3861 -4242
rect 3710 -7907 3861 -7895
rect 3596 -8357 3743 -8345
rect 3269 -8469 3409 -8459
rect 3257 -8524 3269 -8478
rect 3409 -8484 3457 -8478
rect 3445 -8518 3457 -8484
rect 3409 -8524 3457 -8518
rect 3269 -8543 3409 -8533
rect 3170 -8714 3176 -8546
rect 3210 -8571 3216 -8546
rect 3498 -8546 3544 -8534
rect 3498 -8571 3504 -8546
rect 3210 -8689 3504 -8571
rect 3210 -8714 3216 -8689
rect 3170 -8804 3216 -8714
rect 3498 -8714 3504 -8689
rect 3538 -8714 3544 -8546
rect 3305 -8733 3445 -8723
rect 3498 -8726 3544 -8714
rect 3257 -8742 3305 -8736
rect 3257 -8776 3269 -8742
rect 3257 -8782 3305 -8776
rect 3445 -8782 3457 -8736
rect 3305 -8795 3445 -8785
rect 3170 -8972 3176 -8804
rect 3210 -8823 3216 -8804
rect 3498 -8804 3544 -8792
rect 3498 -8823 3504 -8804
rect 3210 -8941 3504 -8823
rect 3210 -8972 3216 -8941
rect 1720 -9063 2763 -9059
rect 1708 -9069 2775 -9063
rect 1708 -9177 1720 -9069
rect 2763 -9177 2775 -9069
rect 1708 -9183 2775 -9177
rect 1720 -9187 2763 -9183
rect 3170 -9203 3216 -8972
rect 3498 -8972 3504 -8941
rect 3538 -8972 3544 -8804
rect 3269 -8985 3409 -8975
rect 3498 -8984 3544 -8972
rect 3257 -9040 3269 -8994
rect 3409 -9000 3457 -8994
rect 3445 -9034 3457 -9000
rect 3409 -9040 3457 -9034
rect 3269 -9059 3409 -9049
rect 3170 -9209 3357 -9203
rect 3170 -9243 3269 -9209
rect 3345 -9243 3357 -9209
rect 3170 -9249 3357 -9243
rect 3170 -9267 3216 -9249
rect 3149 -9271 3216 -9267
rect 3149 -9277 3176 -9271
rect 3210 -9277 3216 -9271
rect 2724 -9302 2884 -9290
rect 1961 -9370 2571 -9332
rect 1961 -9444 1966 -9370
rect 2566 -9444 2571 -9370
rect 1961 -9477 2571 -9444
rect 1961 -9511 2006 -9477
rect 2040 -9511 2106 -9477
rect 2140 -9511 2206 -9477
rect 2240 -9511 2306 -9477
rect 2340 -9511 2406 -9477
rect 2440 -9511 2506 -9477
rect 2540 -9511 2571 -9477
rect 1374 -10083 1498 -10070
rect 1535 -9551 1643 -9539
rect 1535 -10078 1541 -9551
rect 1637 -10078 1643 -9551
rect 1535 -10090 1643 -10078
rect 1961 -9577 2571 -9511
rect 1961 -9611 2006 -9577
rect 2040 -9611 2106 -9577
rect 2140 -9611 2206 -9577
rect 2240 -9611 2306 -9577
rect 2340 -9611 2406 -9577
rect 2440 -9611 2506 -9577
rect 2540 -9611 2571 -9577
rect 1961 -9677 2571 -9611
rect 1961 -9711 2006 -9677
rect 2040 -9711 2106 -9677
rect 2140 -9711 2206 -9677
rect 2240 -9711 2306 -9677
rect 2340 -9711 2406 -9677
rect 2440 -9711 2506 -9677
rect 2540 -9711 2571 -9677
rect 1961 -9777 2571 -9711
rect 1961 -9811 2006 -9777
rect 2040 -9811 2106 -9777
rect 2140 -9811 2206 -9777
rect 2240 -9811 2306 -9777
rect 2340 -9811 2406 -9777
rect 2440 -9811 2506 -9777
rect 2540 -9811 2571 -9777
rect 1961 -9877 2571 -9811
rect 1961 -9911 2006 -9877
rect 2040 -9911 2106 -9877
rect 2140 -9911 2206 -9877
rect 2240 -9911 2306 -9877
rect 2340 -9911 2406 -9877
rect 2440 -9911 2506 -9877
rect 2540 -9911 2571 -9877
rect 1961 -9942 2571 -9911
rect 1961 -10124 2013 -9942
rect 2153 -10098 2632 -10094
rect -93 -10176 2013 -10124
rect 2141 -10104 2644 -10098
rect -1305 -10200 -1153 -10196
rect -315 -10200 -167 -10196
rect -1567 -10275 -1381 -10263
rect -1317 -10206 -1141 -10200
rect -1317 -10260 -1305 -10206
rect -1153 -10260 -1141 -10206
rect -1317 -10266 -1141 -10260
rect -327 -10206 -155 -10200
rect -327 -10260 -315 -10206
rect -167 -10260 -155 -10206
rect 2141 -10224 2153 -10104
rect 2632 -10224 2644 -10104
rect 2724 -10127 2730 -9302
rect 2878 -10127 2884 -9302
rect 3214 -9321 3216 -9277
rect 3398 -9271 3444 -9259
rect 3398 -9321 3404 -9271
rect 3214 -9603 3404 -9321
rect 3214 -9636 3216 -9603
rect 3149 -9639 3176 -9636
rect 3210 -9639 3216 -9636
rect 3149 -9646 3216 -9639
rect 3170 -9721 3216 -9646
rect 3398 -9639 3404 -9603
rect 3438 -9639 3444 -9271
rect 3596 -9343 3602 -8357
rect 3737 -9343 3743 -8357
rect 3596 -9355 3604 -9343
rect 3269 -9658 3345 -9648
rect 3398 -9651 3444 -9639
rect 3257 -9707 3269 -9661
rect 3345 -9707 3357 -9661
rect 3269 -9720 3345 -9710
rect 3149 -9729 3216 -9721
rect 3149 -9731 3176 -9729
rect 3210 -9731 3216 -9729
rect 3214 -9768 3216 -9731
rect 3398 -9729 3444 -9717
rect 3398 -9768 3404 -9729
rect 3214 -10050 3404 -9768
rect 3214 -10090 3216 -10050
rect 3149 -10097 3176 -10090
rect 3210 -10097 3216 -10090
rect 3149 -10100 3216 -10097
rect 2724 -10139 2884 -10127
rect 3170 -10119 3216 -10100
rect 3398 -10097 3404 -10050
rect 3438 -10097 3444 -9729
rect 3398 -10109 3444 -10097
rect 3170 -10125 3357 -10119
rect 3170 -10159 3269 -10125
rect 3345 -10159 3357 -10125
rect 3170 -10165 3357 -10159
rect 2141 -10230 2644 -10224
rect 2153 -10234 2632 -10230
rect -327 -10266 -155 -10260
rect -1305 -10270 -1153 -10266
rect -315 -10270 -167 -10266
rect 3598 -10336 3604 -9355
rect 3736 -9355 3743 -9343
rect 3809 -8356 3969 -8344
rect 3736 -10336 3742 -9355
rect 3598 -10348 3742 -10336
rect 3809 -10335 3815 -8356
rect 3963 -10335 3969 -8356
rect 3809 -10347 3969 -10335
<< via1 >>
rect -1814 7424 778 7627
rect -10213 5416 -2415 5505
rect -6300 4719 -6290 5055
rect -6290 4719 -6256 5055
rect -6256 4719 -6246 5055
rect -9981 4231 -9948 4536
rect -9948 4231 -9914 4536
rect -9914 4231 -9905 4536
rect -6300 4231 -6290 4567
rect -6290 4231 -6256 4567
rect -6256 4231 -6246 4567
rect -2640 4231 -2632 4526
rect -2632 4231 -2598 4526
rect -2598 4231 -2564 4526
rect -1814 4016 -1649 7424
rect -1492 4155 -1476 5155
rect -1476 4155 -1442 5155
rect -1442 4155 -1428 5155
rect -1057 6531 -1038 7131
rect -1038 6531 -1004 7131
rect -1004 6531 -985 7131
rect -615 5392 -600 6392
rect -600 5392 -566 6392
rect -566 5392 -551 6392
rect -181 6531 -162 7131
rect -162 6531 -128 7131
rect -128 6531 -109 7131
rect 261 4155 276 5155
rect 276 4155 310 5155
rect 310 4155 325 5155
rect -1414 4096 -1134 4105
rect -1414 4062 -1134 4096
rect -1414 4053 -1134 4062
rect -976 4096 -696 4105
rect -976 4062 -696 4096
rect -976 4053 -696 4062
rect -538 4096 -258 4105
rect -538 4062 -258 4096
rect -538 4053 -258 4062
rect -100 4096 180 4105
rect -100 4062 180 4096
rect -100 4053 180 4062
rect -9981 3769 -9672 3853
rect -9173 3778 -8824 3845
rect -4109 3775 -3760 3842
rect -1414 3760 -1314 3860
rect -728 3760 -628 3860
rect -290 3760 -190 3860
rect -100 3760 0 3860
rect 1725 3760 2007 3860
rect -8746 3588 -8397 3655
rect -3689 3592 -3340 3659
rect -2975 3589 -2585 3659
rect -1166 3451 -1066 3551
rect -976 3451 -876 3551
rect -538 3451 -438 3551
rect 148 3451 248 3551
rect -1346 3247 -1066 3256
rect -8782 2615 -8738 3183
rect -8738 2615 -8704 3183
rect -8704 2615 -8696 3183
rect -6288 2039 -6280 2358
rect -6280 2039 -6246 2358
rect -6246 2039 -6236 2358
rect -1346 3213 -1066 3247
rect -1346 3204 -1066 3213
rect -908 3247 -628 3256
rect -908 3213 -628 3247
rect -908 3204 -628 3213
rect -470 3247 -190 3256
rect -470 3213 -190 3247
rect -470 3204 -190 3213
rect -32 3247 248 3256
rect -32 3213 248 3247
rect -32 3204 248 3213
rect -3830 2615 -3822 3183
rect -3822 2615 -3788 3183
rect -3788 2615 -3744 3183
rect -8672 1957 -8462 1969
rect -8672 1923 -8462 1957
rect -8672 1912 -8462 1923
rect -4060 1957 -3850 1969
rect -4060 1923 -3850 1957
rect -4060 1912 -3850 1923
rect -8649 1794 -8462 1851
rect -6219 1791 -6018 1855
rect -10065 1670 -9489 1687
rect -10065 1636 -9489 1670
rect -10065 1632 -9489 1636
rect -6519 1479 -6309 1536
rect -4060 1481 -3850 1538
rect -9447 640 -9439 1439
rect -9439 640 -9405 1439
rect -9405 640 -9395 1439
rect -6519 1392 -6309 1404
rect -6519 1358 -6309 1392
rect -6519 1347 -6309 1358
rect -6219 1392 -6009 1403
rect -6219 1358 -6009 1392
rect -8849 236 -8739 1308
rect -8739 236 -8705 1308
rect -8705 236 -8697 1308
rect -6219 1346 -6009 1358
rect -6289 958 -6281 1277
rect -6281 958 -6247 1277
rect -6247 958 -6237 1277
rect -10291 -26 -9738 68
rect -8677 82 -8197 89
rect -8677 48 -8197 82
rect -8677 37 -8197 48
rect -6219 82 -5739 90
rect -3832 236 -3823 1308
rect -3823 236 -3789 1308
rect -3789 236 -3680 1308
rect -6219 48 -5739 82
rect -6219 38 -5739 48
rect -1797 22 -1649 3198
rect -1798 -11 -1649 22
rect -1491 2154 -1476 3154
rect -1476 2154 -1442 3154
rect -1442 2154 -1427 3154
rect -1057 178 -1038 778
rect -1038 178 -1004 778
rect -1004 178 -985 778
rect -615 994 -600 1994
rect -600 994 -566 1994
rect -566 994 -551 1994
rect -182 178 -162 778
rect -162 178 -128 778
rect -128 178 -110 778
rect 261 2154 276 3154
rect 276 2154 310 3154
rect 310 2154 325 3154
rect 11789 2772 12048 2773
rect 7086 2408 12048 2772
rect 7086 2407 11890 2408
rect 1861 1822 5524 2113
rect -1798 -154 767 -11
rect -1685 -155 767 -154
rect -10289 -256 -3355 -167
rect 3344 600 3353 1600
rect 3353 600 3387 1600
rect 3387 600 3396 1600
rect 3762 224 3771 1224
rect 3771 224 3805 1224
rect 3805 224 3814 1224
rect 4180 600 4189 1600
rect 4189 600 4223 1600
rect 4223 600 4232 1600
rect 4598 224 4607 1224
rect 4607 224 4641 1224
rect 4641 224 4650 1224
rect 5016 600 5025 1600
rect 5025 600 5059 1600
rect 5059 600 5068 1600
rect 5237 306 5524 1822
rect 5224 121 5348 180
rect 7148 205 7265 2407
rect 7431 1669 7446 1869
rect 7446 1669 7480 1869
rect 7480 1669 7495 1869
rect 8495 1845 8504 2145
rect 8504 1845 8538 2145
rect 8538 1845 8547 2145
rect 9547 1945 9562 2145
rect 9562 1945 9596 2145
rect 9596 1945 9611 2145
rect 10611 1845 10620 2145
rect 10620 1845 10654 2145
rect 10654 1845 10663 2145
rect 11663 1669 11678 1869
rect 11678 1669 11712 1869
rect 11712 1669 11727 1869
rect 7836 1610 8476 1619
rect 7836 1576 8476 1610
rect 7836 1567 8476 1576
rect 8894 1610 9534 1619
rect 9952 1610 10592 1620
rect 8894 1576 9534 1610
rect 9952 1576 10592 1610
rect 8894 1567 9534 1576
rect 9952 1568 10592 1576
rect 11010 1610 11650 1619
rect 11010 1576 11650 1610
rect 11010 1567 11650 1576
rect 11932 1594 12029 2408
rect 8376 1371 8476 1471
rect 8566 1371 8666 1471
rect 9624 1371 9724 1471
rect 11550 1371 11650 1471
rect 7508 1189 7608 1289
rect 9434 1189 9534 1289
rect 10492 1189 10592 1289
rect 10682 1189 10782 1289
rect 7508 1076 8148 1085
rect 7508 1042 8148 1076
rect 7508 1033 8148 1042
rect 8566 1076 9206 1085
rect 9624 1076 10264 1085
rect 8566 1042 9206 1076
rect 9624 1042 10264 1076
rect 8566 1033 9206 1042
rect 9624 1033 10264 1042
rect 10682 1076 11322 1085
rect 10682 1042 11322 1076
rect 10682 1033 11322 1042
rect 7431 783 7446 983
rect 7446 783 7480 983
rect 7480 783 7495 983
rect 8495 507 8504 807
rect 8504 507 8538 807
rect 8538 507 8547 807
rect 9547 507 9562 707
rect 9562 507 9596 707
rect 9596 507 9611 707
rect 10611 507 10620 807
rect 10620 507 10654 807
rect 10654 507 10663 807
rect 11663 783 11678 983
rect 11678 783 11712 983
rect 11712 783 11727 983
rect 7148 115 11697 205
rect 7183 108 11697 115
rect 3071 -170 5134 66
rect -1742 -501 -1595 -493
rect -1742 -502 -1466 -501
rect 6078 -502 6084 -456
rect 6084 -502 6200 -456
rect -1742 -605 6200 -502
rect -1742 -1795 -1595 -605
rect 6078 -617 6084 -605
rect 6084 -617 6200 -605
rect 6200 -617 6225 -456
rect 6078 -639 6225 -617
rect 8506 -128 10634 -25
rect 8506 -666 8564 -128
rect 9080 -462 9089 -302
rect 9089 -462 9123 -302
rect 9123 -462 9132 -302
rect -1481 -972 -1466 -872
rect -1466 -972 -1432 -872
rect -1432 -972 -1417 -872
rect 463 -972 472 -872
rect 472 -972 506 -872
rect 506 -972 515 -872
rect 2395 -1148 2410 -1048
rect 2410 -1148 2444 -1048
rect 2444 -1148 2459 -1048
rect 4339 -972 4348 -872
rect 4348 -972 4382 -872
rect 4382 -972 4391 -872
rect 8599 -868 8631 -731
rect 8631 -868 8665 -731
rect 8665 -868 8693 -731
rect 6271 -972 6286 -872
rect 6286 -972 6320 -872
rect 6320 -972 6335 -872
rect 9996 -462 10005 -302
rect 10005 -462 10039 -302
rect 10039 -462 10048 -302
rect 9518 -610 9547 -473
rect 9547 -610 9581 -473
rect 9581 -610 9612 -473
rect 10434 -868 10463 -731
rect 10463 -868 10497 -731
rect 10497 -868 10528 -731
rect 8861 -928 9061 -919
rect 8861 -962 9061 -928
rect 8861 -971 9061 -962
rect 9319 -928 9519 -919
rect 9319 -962 9519 -928
rect 9319 -971 9519 -962
rect 9777 -928 9977 -919
rect 9777 -962 9977 -928
rect 9777 -971 9977 -962
rect 10235 -928 10435 -919
rect 10235 -962 10435 -928
rect 10235 -971 10435 -962
rect 7122 -1143 7205 -1043
rect 8961 -1143 9061 -1043
rect 9151 -1143 9251 -1043
rect 9609 -1143 9709 -1043
rect 10335 -1143 10435 -1043
rect -1481 -1558 -1466 -1458
rect -1466 -1558 -1432 -1458
rect -1432 -1558 -1417 -1458
rect 463 -1558 472 -1458
rect 472 -1558 506 -1458
rect 506 -1558 515 -1458
rect 2395 -1382 2410 -1282
rect 2410 -1382 2444 -1282
rect 2444 -1382 2459 -1282
rect 4339 -1558 4348 -1458
rect 4348 -1558 4382 -1458
rect 4382 -1558 4391 -1458
rect 7112 -1329 7225 -1229
rect 8693 -1329 8793 -1229
rect 9419 -1329 9519 -1229
rect 9877 -1329 9977 -1229
rect 10067 -1329 10167 -1229
rect 6271 -1558 6286 -1458
rect 6286 -1558 6320 -1458
rect 6320 -1558 6335 -1458
rect 8693 -1425 8893 -1416
rect 8693 -1459 8893 -1425
rect 8693 -1468 8893 -1459
rect 9151 -1425 9351 -1416
rect 9151 -1459 9351 -1425
rect 9151 -1468 9351 -1459
rect 9609 -1425 9809 -1416
rect 9609 -1459 9809 -1425
rect 9609 -1468 9809 -1459
rect 10067 -1425 10267 -1416
rect 10067 -1459 10267 -1425
rect 10067 -1468 10267 -1459
rect 8600 -1657 8631 -1520
rect 8631 -1657 8665 -1520
rect 8665 -1657 8694 -1520
rect -1742 -1796 -1501 -1795
rect -1742 -1993 6177 -1796
rect 8497 -2333 8571 -1702
rect 9517 -1868 9547 -1731
rect 9547 -1868 9581 -1731
rect 9581 -1868 9611 -1731
rect 9080 -2085 9089 -1925
rect 9089 -2085 9123 -1925
rect 9123 -2085 9132 -1925
rect 10432 -1657 10463 -1520
rect 10463 -1657 10497 -1520
rect 10497 -1657 10526 -1520
rect 9996 -2085 10005 -1925
rect 10005 -2085 10039 -1925
rect 10039 -2085 10048 -1925
rect 11593 -1051 11697 108
rect 11770 -620 11779 -420
rect 11779 -620 11813 -420
rect 11813 -620 11822 -420
rect 12126 -620 12135 -420
rect 12135 -620 12169 -420
rect 12169 -620 12178 -420
rect 11898 -916 11907 -716
rect 11907 -916 11941 -716
rect 11941 -916 11950 -716
rect 12254 -916 12263 -716
rect 12263 -916 12297 -716
rect 12297 -916 12306 -716
rect 11898 -1381 11950 -1302
rect 11810 -1601 11819 -1530
rect 11819 -1601 11853 -1530
rect 11853 -1601 11862 -1530
rect 12254 -1496 12263 -1425
rect 12263 -1496 12297 -1425
rect 12297 -1496 12306 -1425
rect 12166 -1601 12175 -1530
rect 12175 -1601 12209 -1530
rect 12209 -1601 12218 -1530
rect 10997 -2157 12375 -1885
rect 3710 -2900 3861 -2888
rect -1561 -10263 -1387 -3685
rect -1136 -3815 -936 -3800
rect -1136 -3849 -936 -3815
rect 921 -3815 1121 -3806
rect -1136 -3864 -936 -3849
rect -319 -3977 -310 -3877
rect -310 -3977 -276 -3877
rect -276 -3977 -267 -3877
rect -93 -3929 -41 -3829
rect -560 -4073 -360 -4062
rect -560 -4107 -360 -4073
rect -560 -4118 -360 -4107
rect -93 -4187 -41 -4087
rect -784 -4331 -684 -4322
rect -784 -4365 -684 -4331
rect -784 -4374 -684 -4365
rect -790 -4503 -685 -4451
rect -319 -4493 -310 -4393
rect -310 -4493 -276 -4393
rect -276 -4493 -267 -4393
rect -1136 -4589 -936 -4580
rect -1136 -4623 -936 -4589
rect -1136 -4632 -936 -4623
rect -787 -4765 -687 -4713
rect -784 -4847 -684 -4838
rect -784 -4881 -684 -4847
rect -784 -4890 -684 -4881
rect -319 -5034 -310 -4909
rect -310 -5034 -276 -4909
rect -276 -5034 -267 -4909
rect -93 -4961 -41 -4861
rect -560 -5105 -360 -5094
rect -560 -5139 -360 -5105
rect -560 -5150 -360 -5139
rect -1136 -5363 -936 -5348
rect -1136 -5397 -936 -5363
rect -1136 -5412 -936 -5397
rect -560 -5621 -360 -5610
rect -560 -5655 -360 -5621
rect -560 -5666 -360 -5655
rect -93 -5735 -41 -5635
rect -784 -5879 -684 -5870
rect -784 -5913 -684 -5879
rect -784 -5922 -684 -5913
rect -785 -6056 -685 -6004
rect -319 -6041 -310 -5941
rect -310 -6041 -276 -5941
rect -276 -6041 -267 -5941
rect -1136 -6137 -936 -6129
rect -1136 -6171 -936 -6137
rect -1136 -6181 -936 -6171
rect -782 -6308 -682 -6256
rect -784 -6395 -684 -6386
rect -784 -6429 -684 -6395
rect -784 -6438 -684 -6429
rect -319 -6583 -310 -6457
rect -310 -6583 -276 -6457
rect -276 -6583 -267 -6457
rect -93 -6509 -41 -6409
rect -560 -6653 -360 -6642
rect -560 -6687 -360 -6653
rect -560 -6698 -360 -6687
rect -1136 -6911 -936 -6896
rect -1136 -6945 -936 -6911
rect -1136 -6960 -936 -6945
rect -560 -7169 -360 -7158
rect -560 -7203 -360 -7169
rect -560 -7214 -360 -7203
rect -93 -7283 -41 -7183
rect -784 -7427 -684 -7418
rect -784 -7461 -684 -7427
rect -784 -7470 -684 -7461
rect -783 -7601 -683 -7549
rect -319 -7589 -310 -7489
rect -310 -7589 -276 -7489
rect -276 -7589 -267 -7489
rect -1136 -7685 -936 -7676
rect -1136 -7719 -936 -7685
rect -1136 -7728 -936 -7719
rect -785 -7863 -685 -7811
rect -784 -7943 -684 -7934
rect -784 -7977 -684 -7943
rect -784 -7986 -684 -7977
rect -319 -8131 -310 -8005
rect -310 -8131 -276 -8005
rect -276 -8131 -267 -8005
rect -93 -8057 -41 -7957
rect -560 -8201 -360 -8190
rect -560 -8235 -360 -8201
rect -560 -8246 -360 -8235
rect -1136 -8459 -936 -8444
rect -1136 -8493 -936 -8459
rect -1136 -8508 -936 -8493
rect -560 -8717 -360 -8706
rect -560 -8751 -360 -8717
rect -560 -8762 -360 -8751
rect -93 -8831 -41 -8731
rect -784 -8975 -684 -8966
rect -784 -9009 -684 -8975
rect -784 -9018 -684 -9009
rect -784 -9145 -684 -9093
rect -319 -9137 -310 -9037
rect -310 -9137 -276 -9037
rect -276 -9137 -267 -9037
rect -1136 -9233 -936 -9224
rect -1136 -9267 -936 -9233
rect -1136 -9276 -936 -9267
rect -784 -9410 -684 -9358
rect -784 -9491 -684 -9482
rect -784 -9525 -684 -9491
rect -784 -9534 -684 -9525
rect -319 -9653 -310 -9553
rect -310 -9653 -276 -9553
rect -276 -9653 -267 -9553
rect -93 -9605 -41 -9505
rect -560 -9749 -360 -9738
rect -560 -9783 -360 -9749
rect -560 -9794 -360 -9783
rect -1136 -10007 -936 -9992
rect -1136 -10041 -936 -10007
rect -1136 -10056 -936 -10041
rect 52 -3929 104 -3829
rect 921 -3849 1121 -3815
rect 921 -3858 1121 -3849
rect 252 -3977 261 -3877
rect 261 -3977 295 -3877
rect 295 -3977 304 -3877
rect 644 -3990 744 -3938
rect 646 -4073 746 -4064
rect 646 -4107 746 -4073
rect 646 -4116 746 -4107
rect 252 -4303 261 -4135
rect 261 -4303 295 -4135
rect 295 -4303 304 -4135
rect 252 -4319 304 -4303
rect 52 -4445 104 -4345
rect 921 -4331 1121 -4320
rect 921 -4365 1121 -4331
rect 921 -4376 1121 -4365
rect 345 -4589 545 -4574
rect 345 -4623 545 -4589
rect 345 -4638 545 -4623
rect 921 -4847 1121 -4836
rect 921 -4881 1121 -4847
rect 921 -4892 1121 -4881
rect 52 -5219 104 -5119
rect 646 -5105 746 -5096
rect 646 -5139 746 -5105
rect 646 -5148 746 -5139
rect 252 -5267 261 -5167
rect 261 -5267 295 -5167
rect 295 -5267 304 -5167
rect 646 -5282 746 -5230
rect 921 -5363 1121 -5354
rect 921 -5397 1121 -5363
rect 921 -5406 1121 -5397
rect 648 -5537 748 -5485
rect 646 -5621 746 -5612
rect 646 -5655 746 -5621
rect 646 -5664 746 -5655
rect 252 -5851 261 -5683
rect 261 -5851 295 -5683
rect 295 -5851 304 -5683
rect 252 -5867 304 -5851
rect 52 -5993 104 -5893
rect 921 -5879 1121 -5868
rect 921 -5913 1121 -5879
rect 921 -5924 1121 -5913
rect 345 -6137 545 -6122
rect 345 -6171 545 -6137
rect 345 -6186 545 -6171
rect 921 -6395 1121 -6384
rect 921 -6429 1121 -6395
rect 921 -6440 1121 -6429
rect 52 -6767 104 -6667
rect 645 -6653 745 -6644
rect 645 -6687 745 -6653
rect 645 -6696 745 -6687
rect 252 -6815 261 -6715
rect 261 -6815 295 -6715
rect 295 -6815 304 -6715
rect 648 -6833 748 -6781
rect 921 -6911 1121 -6902
rect 921 -6945 1121 -6911
rect 921 -6954 1121 -6945
rect 646 -7095 746 -7043
rect 646 -7169 746 -7160
rect 646 -7203 746 -7169
rect 646 -7212 746 -7203
rect 252 -7399 261 -7231
rect 261 -7399 295 -7231
rect 295 -7399 304 -7231
rect 252 -7415 304 -7399
rect 52 -7541 104 -7441
rect 921 -7427 1121 -7416
rect 921 -7461 1121 -7427
rect 921 -7472 1121 -7461
rect 345 -7685 545 -7670
rect 345 -7719 545 -7685
rect 345 -7734 545 -7719
rect 921 -7943 1121 -7932
rect 921 -7977 1121 -7943
rect 921 -7988 1121 -7977
rect 52 -8315 104 -8215
rect 646 -8201 746 -8192
rect 646 -8235 746 -8201
rect 646 -8244 746 -8235
rect 252 -8363 261 -8263
rect 261 -8363 295 -8263
rect 295 -8363 304 -8263
rect 644 -8381 744 -8329
rect 921 -8459 1121 -8450
rect 921 -8493 1121 -8459
rect 921 -8502 1121 -8493
rect 645 -8637 745 -8585
rect 646 -8717 746 -8708
rect 646 -8751 746 -8717
rect 646 -8760 746 -8751
rect 252 -8947 261 -8779
rect 261 -8947 295 -8779
rect 295 -8947 304 -8779
rect 252 -8979 304 -8947
rect 921 -8975 1121 -8964
rect 52 -9089 104 -8989
rect 921 -9009 1121 -8975
rect 921 -9020 1121 -9009
rect 345 -9233 545 -9218
rect 345 -9267 545 -9233
rect 345 -9282 545 -9267
rect 920 -9491 1120 -9480
rect 920 -9525 1120 -9491
rect 920 -9536 1120 -9525
rect 52 -9863 104 -9763
rect 646 -9749 746 -9740
rect 646 -9783 746 -9749
rect 646 -9792 746 -9783
rect 252 -9911 261 -9811
rect 261 -9911 295 -9811
rect 295 -9911 304 -9811
rect 648 -9915 748 -9863
rect 921 -10007 1121 -9998
rect 921 -10041 1121 -10007
rect 921 -10050 1121 -10041
rect 1380 -10070 1492 -3729
rect 2122 -8325 2313 -2918
rect 3269 -2945 3392 -2936
rect 3269 -2979 3392 -2945
rect 3269 -2988 3392 -2979
rect 2482 -3010 2542 -3001
rect 2598 -3010 2658 -3001
rect 2482 -3044 2542 -3010
rect 2598 -3044 2658 -3010
rect 2482 -3053 2542 -3044
rect 2598 -3053 2658 -3044
rect 2598 -3268 2658 -3259
rect 2598 -3302 2658 -3268
rect 2598 -3311 2658 -3302
rect 2482 -3526 2542 -3517
rect 2482 -3560 2542 -3526
rect 2482 -3569 2542 -3560
rect 2598 -3784 2658 -3775
rect 2598 -3818 2658 -3784
rect 2598 -3827 2658 -3818
rect 2482 -4042 2542 -4033
rect 2482 -4076 2542 -4042
rect 2482 -4085 2542 -4076
rect 3322 -3403 3445 -3394
rect 3322 -3437 3445 -3403
rect 3322 -3446 3445 -3437
rect 3269 -3526 3392 -3517
rect 3269 -3560 3392 -3526
rect 3269 -3569 3392 -3560
rect 2482 -4300 2542 -4291
rect 2482 -4334 2542 -4300
rect 2482 -4343 2542 -4334
rect 2598 -4558 2658 -4549
rect 2598 -4592 2658 -4558
rect 2598 -4601 2658 -4592
rect 2482 -4816 2542 -4807
rect 2482 -4850 2542 -4816
rect 2482 -4859 2542 -4850
rect 2598 -5074 2658 -5065
rect 2598 -5108 2658 -5074
rect 2598 -5117 2658 -5108
rect 2482 -5332 2542 -5323
rect 2482 -5366 2542 -5332
rect 2482 -5375 2542 -5366
rect 3321 -3984 3445 -3975
rect 3321 -4018 3445 -3984
rect 3321 -4027 3445 -4018
rect 3710 -4242 3716 -2900
rect 3269 -4816 3382 -4807
rect 3269 -4850 3382 -4816
rect 3269 -4859 3382 -4850
rect 2482 -5590 2542 -5581
rect 2482 -5624 2542 -5590
rect 2482 -5633 2542 -5624
rect 2598 -5848 2658 -5839
rect 2598 -5882 2658 -5848
rect 2598 -5891 2658 -5882
rect 2482 -6106 2542 -6097
rect 2482 -6140 2542 -6106
rect 2482 -6149 2542 -6140
rect 2598 -6364 2658 -6355
rect 2598 -6398 2658 -6364
rect 2598 -6407 2658 -6398
rect 2482 -6622 2542 -6613
rect 2482 -6656 2542 -6622
rect 2482 -6665 2542 -6656
rect 3322 -5274 3445 -5265
rect 3322 -5308 3445 -5274
rect 3322 -5317 3445 -5308
rect 3269 -6106 3382 -6097
rect 3269 -6140 3382 -6106
rect 3269 -6149 3382 -6140
rect 2482 -6880 2542 -6871
rect 2482 -6914 2542 -6880
rect 2482 -6923 2542 -6914
rect 2598 -7138 2658 -7129
rect 2598 -7172 2658 -7138
rect 2598 -7181 2658 -7172
rect 2482 -7396 2542 -7387
rect 2482 -7430 2542 -7396
rect 2482 -7439 2542 -7430
rect 2598 -7654 2658 -7645
rect 2598 -7688 2658 -7654
rect 2598 -7697 2658 -7688
rect 2482 -7912 2542 -7903
rect 2482 -7946 2542 -7912
rect 2482 -7955 2542 -7946
rect 3322 -6564 3445 -6555
rect 3322 -6598 3445 -6564
rect 3322 -6607 3445 -6598
rect 3269 -7396 3382 -7387
rect 3269 -7430 3382 -7396
rect 3269 -7439 3382 -7430
rect 2482 -8170 2542 -8161
rect 2482 -8204 2542 -8170
rect 2482 -8213 2542 -8204
rect 3322 -7854 3445 -7845
rect 3322 -7888 3445 -7854
rect 3322 -7897 3445 -7888
rect 3716 -7895 3855 -2900
rect 3855 -4242 3861 -2900
rect 8452 -2340 8679 -2333
rect 8452 -2503 9795 -2340
rect 8452 -3519 8790 -2503
rect 8790 -2510 9795 -2503
rect 9719 -2635 10128 -2619
rect 9719 -2669 10128 -2635
rect 9719 -2684 10128 -2669
rect 8957 -2852 8968 -2712
rect 8968 -2852 9002 -2712
rect 9002 -2852 9013 -2712
rect 9052 -2993 9552 -2978
rect 9052 -3027 9552 -2993
rect 9052 -3042 9552 -3027
rect 9719 -3351 10128 -3335
rect 9719 -3385 10128 -3351
rect 9719 -3400 10128 -3385
rect 10341 -3519 10552 -2468
rect 11293 -2385 11495 -2377
rect 11293 -2423 11495 -2385
rect 11293 -2429 11495 -2423
rect 12127 -2385 12329 -2378
rect 12127 -2423 12329 -2385
rect 12127 -2430 12329 -2423
rect 8452 -3758 10552 -3519
rect 8452 -3760 8679 -3758
rect 10341 -3769 10552 -3758
rect 3269 -8484 3409 -8469
rect 3269 -8518 3409 -8484
rect 3269 -8533 3409 -8518
rect 3305 -8742 3445 -8733
rect 3305 -8776 3445 -8742
rect 3305 -8785 3445 -8776
rect 1720 -9177 2763 -9069
rect 3269 -9000 3409 -8985
rect 3269 -9034 3409 -9000
rect 3269 -9049 3409 -9034
rect 1966 -9377 2566 -9370
rect 1966 -9411 2006 -9377
rect 2006 -9411 2040 -9377
rect 2040 -9411 2106 -9377
rect 2106 -9411 2140 -9377
rect 2140 -9411 2206 -9377
rect 2206 -9411 2240 -9377
rect 2240 -9411 2306 -9377
rect 2306 -9411 2340 -9377
rect 2340 -9411 2406 -9377
rect 2406 -9411 2440 -9377
rect 2440 -9411 2506 -9377
rect 2506 -9411 2540 -9377
rect 2540 -9411 2566 -9377
rect 1966 -9444 2566 -9411
rect 1541 -10078 1637 -9551
rect -1305 -10260 -1153 -10206
rect -315 -10260 -167 -10206
rect 2153 -10224 2632 -10104
rect 2730 -10127 2878 -9302
rect 3149 -9636 3176 -9277
rect 3176 -9636 3210 -9277
rect 3210 -9636 3214 -9277
rect 3602 -8444 3637 -8357
rect 3637 -8444 3737 -8357
rect 3602 -9343 3737 -8444
rect 3269 -9667 3345 -9658
rect 3269 -9701 3345 -9667
rect 3269 -9710 3345 -9701
rect 3149 -10090 3176 -9731
rect 3176 -10090 3210 -9731
rect 3210 -10090 3214 -9731
rect 3604 -10336 3736 -9343
rect 3815 -10335 3963 -8356
<< metal2 >>
rect -1903 7627 778 7637
rect -1903 7413 -1814 7627
rect -2376 5806 -1814 5808
rect -10397 5505 -1814 5806
rect -10397 5416 -10213 5505
rect -2415 5416 -1814 5505
rect -10397 5406 -1814 5416
rect -6300 5055 -6246 5406
rect -2376 5405 -1814 5406
rect -9991 4536 -9905 4579
rect -9991 4231 -9981 4536
rect -9991 3863 -9905 4231
rect -6300 4567 -6246 4719
rect -6300 4221 -6246 4231
rect -2640 4526 -2554 4579
rect -2564 4231 -2554 4526
rect -9991 3853 -9672 3863
rect -9991 3769 -9981 3853
rect -9991 3759 -9672 3769
rect -9173 3845 -8812 3860
rect -8824 3778 -8812 3845
rect -9173 3760 -8812 3778
rect -4109 3842 -3744 3860
rect -3760 3775 -3744 3842
rect -4109 3760 -3744 3775
rect -10065 1697 -9489 1707
rect -10065 1622 -9489 1632
rect -9447 1448 -9395 1449
rect -9450 1439 -9392 1448
rect -9450 1438 -9447 1439
rect -9395 1438 -9392 1439
rect -9450 630 -9392 640
rect -8898 1318 -8812 3760
rect -8782 3655 -8396 3675
rect -8782 3588 -8746 3655
rect -8397 3588 -8396 3655
rect -8782 3575 -8396 3588
rect -8782 3183 -8696 3575
rect -8782 2605 -8696 2615
rect -3830 3183 -3744 3760
rect -2640 3675 -2554 4231
rect -1649 7414 778 7424
rect -1057 7131 1624 7141
rect -985 7041 -181 7131
rect -1057 6521 -985 6531
rect -109 7041 1624 7131
rect -181 6521 -109 6531
rect -615 6392 -551 6402
rect -615 5382 -551 5392
rect -1492 5155 -1428 5165
rect -1492 4145 -1428 4155
rect 261 5155 325 5165
rect 261 4145 325 4155
rect -1814 4006 -1649 4016
rect -1414 4105 -1134 4115
rect -1414 4043 -1134 4053
rect -976 4105 -696 4115
rect -976 4043 -696 4053
rect -538 4105 -258 4115
rect -538 4043 -258 4053
rect -100 4105 180 4115
rect -100 4043 180 4053
rect -1414 3860 -1314 4043
rect -1414 3750 -1314 3760
rect -3830 2605 -3744 2615
rect -3714 3659 -3340 3675
rect -3714 3592 -3689 3659
rect -3714 3575 -3340 3592
rect -2975 3659 -2554 3675
rect -2585 3589 -2554 3659
rect -2975 3575 -2554 3589
rect -6292 2371 -6236 2381
rect -6292 2019 -6236 2029
rect -8672 1969 -8462 1979
rect -8672 1851 -8462 1912
rect -4060 1969 -3850 1979
rect -8672 1794 -8649 1851
rect -8672 1784 -8462 1794
rect -6219 1855 -6009 1867
rect -6018 1791 -6009 1855
rect -6519 1536 -6309 1546
rect -6519 1404 -6309 1479
rect -6519 1337 -6309 1347
rect -6219 1403 -6009 1791
rect -4060 1538 -3850 1912
rect -4060 1471 -3850 1481
rect -6219 1336 -6009 1346
rect -3714 1318 -3628 3575
rect -1166 3551 -1066 3561
rect -1166 3266 -1066 3451
rect -976 3551 -876 4043
rect -976 3441 -876 3451
rect -728 3860 -628 3870
rect -728 3266 -628 3760
rect -538 3551 -438 4043
rect -538 3441 -438 3451
rect -290 3860 -190 3870
rect -290 3266 -190 3760
rect -100 3860 0 4043
rect -100 3750 0 3760
rect 148 3551 248 3561
rect 148 3266 248 3451
rect -1346 3256 -1066 3266
rect -8898 1308 -8697 1318
rect -8898 236 -8849 1308
rect -3832 1308 -3628 1318
rect -6293 1287 -6235 1297
rect -6293 938 -6235 948
rect -8697 236 -8695 744
rect -8898 167 -8695 236
rect -3680 236 -3628 1308
rect -3832 226 -3628 236
rect -1797 3198 -1649 3208
rect -10599 134 -10501 144
rect -10501 68 -9617 134
rect -10501 -26 -10291 68
rect -9738 -26 -9617 68
rect -8677 92 -8197 102
rect -8677 24 -8197 34
rect -6219 94 -5739 104
rect -6219 26 -5739 36
rect -10501 -157 -9617 -26
rect -1798 22 -1797 32
rect -1346 3194 -1066 3204
rect -908 3256 -628 3266
rect -908 3194 -628 3204
rect -470 3256 -190 3266
rect -470 3194 -190 3204
rect -32 3256 248 3266
rect -32 3194 248 3204
rect -1491 3154 -1427 3164
rect -1491 2144 -1427 2154
rect 261 3154 325 3164
rect 261 2144 325 2154
rect -615 1994 -551 2004
rect -615 984 -551 994
rect 1524 1610 1624 7041
rect 1715 3860 2007 3870
rect 1715 3750 2007 3760
rect 13414 2786 13712 2796
rect 5125 2782 7137 2786
rect 12075 2784 13414 2785
rect 12028 2783 13414 2784
rect 11789 2782 13414 2783
rect 5125 2773 13414 2782
rect 5125 2772 11789 2773
rect 5125 2407 7086 2772
rect 12048 2408 13414 2773
rect 11890 2407 11932 2408
rect 5125 2396 7148 2407
rect 5125 2123 5524 2396
rect 7078 2368 7148 2396
rect 1861 2113 5524 2123
rect 1861 1812 5237 1822
rect 1524 1600 5068 1610
rect 1524 1510 3344 1600
rect -1057 788 343 789
rect 1524 788 1624 1510
rect -1057 778 1624 788
rect -985 689 -182 778
rect -1057 168 -985 178
rect -110 689 1624 778
rect 215 688 1624 689
rect 3396 1510 4180 1600
rect 3344 590 3396 600
rect 3762 1224 3814 1234
rect -182 168 -110 178
rect 4232 1510 5016 1600
rect 4180 590 4232 600
rect 4598 1224 4650 1234
rect 3762 76 3814 224
rect 5016 590 5068 600
rect 5237 296 5524 306
rect 4598 76 4650 224
rect 7265 2398 11932 2407
rect 7265 2397 11890 2398
rect 7265 2368 7293 2397
rect 8495 2145 8547 2397
rect 7431 1869 7495 1879
rect 9547 2145 9611 2155
rect 9547 1935 9611 1945
rect 10611 2145 10663 2397
rect 8495 1835 8547 1845
rect 10611 1835 10663 1845
rect 11663 1869 11727 1879
rect 7431 1659 7495 1669
rect 11663 1659 11727 1669
rect 7836 1619 8476 1629
rect 7836 1557 8476 1567
rect 8894 1619 9534 1629
rect 8894 1557 9534 1567
rect 9952 1620 10592 1630
rect 9952 1558 10592 1568
rect 8376 1471 8476 1557
rect 8376 1361 8476 1371
rect 8566 1471 8666 1481
rect 7508 1289 7608 1299
rect 7508 1095 7608 1189
rect 8566 1095 8666 1371
rect 9434 1289 9534 1557
rect 9434 1179 9534 1189
rect 9624 1471 9724 1481
rect 9624 1095 9724 1371
rect 10492 1289 10592 1558
rect 11010 1619 11650 1629
rect 12029 2399 13414 2408
rect 12029 2398 12048 2399
rect 13414 2389 13712 2399
rect 11932 1584 12029 1594
rect 11010 1557 11650 1567
rect 11550 1471 11650 1557
rect 11550 1361 11650 1371
rect 10492 1179 10592 1189
rect 10682 1289 10782 1299
rect 10682 1095 10782 1189
rect 7508 1085 8148 1095
rect 7508 1023 8148 1033
rect 8566 1085 9206 1095
rect 8566 1023 9206 1033
rect 9624 1085 10264 1095
rect 9624 1023 10264 1033
rect 10682 1085 11322 1095
rect 10682 1023 11322 1033
rect 7431 983 7495 993
rect 11663 983 11727 993
rect 7431 773 7495 783
rect 8495 807 8547 817
rect 10611 807 10663 817
rect 8495 215 8547 507
rect 9547 707 9611 717
rect 9547 497 9611 507
rect 11663 773 11727 783
rect 10611 215 10663 507
rect 7265 205 11697 215
rect 5224 180 6836 190
rect 5348 121 6836 180
rect 5224 111 6836 121
rect 3071 66 5134 76
rect -1649 -11 767 -1
rect -1798 -155 -1685 -154
rect -10501 -167 -3355 -157
rect -1798 -164 767 -155
rect -1685 -165 767 -164
rect -10501 -256 -10289 -167
rect 3071 -180 5134 -170
rect -10501 -266 -3355 -256
rect -10599 -276 -10501 -266
rect -3764 -490 -3355 -266
rect 6078 -456 6225 -446
rect -1742 -490 -1595 -483
rect -3767 -491 -1595 -490
rect -3767 -492 -1466 -491
rect -3767 -493 6078 -492
rect -3767 -827 -1742 -493
rect -1595 -501 6078 -493
rect -1466 -502 6078 -501
rect -1808 -1993 -1742 -1785
rect -1595 -615 6078 -605
rect -1481 -872 -1417 -862
rect -1481 -982 -1417 -972
rect 463 -872 515 -615
rect 463 -982 515 -972
rect 4339 -872 4391 -615
rect 6078 -649 6225 -639
rect 4339 -982 4391 -972
rect 6271 -872 6335 -862
rect 6271 -982 6335 -972
rect 2395 -1048 2459 -1038
rect 2395 -1158 2459 -1148
rect 2395 -1282 2459 -1272
rect 2395 -1392 2459 -1382
rect -1481 -1458 -1417 -1448
rect -1481 -1568 -1417 -1558
rect 463 -1458 515 -1448
rect -1595 -1786 -1501 -1785
rect 463 -1786 515 -1558
rect 4339 -1458 4391 -1448
rect 4339 -1786 4391 -1558
rect 6271 -1458 6335 -1448
rect 6271 -1568 6335 -1558
rect 6245 -1786 6429 -1776
rect -1595 -1795 6245 -1786
rect -1501 -1796 6245 -1795
rect 6177 -1993 6245 -1796
rect -1808 -2003 6245 -1993
rect 6429 -2003 6438 -1786
rect -1572 -3685 -1377 -2003
rect 6245 -2013 6429 -2003
rect 2962 -2314 3062 -2304
rect 2962 -2707 3062 -2494
rect -1572 -3871 -1561 -3685
rect -1571 -10263 -1561 -3871
rect -1387 -4580 -1377 -3685
rect -794 -3646 756 -3526
rect -1146 -3864 -1136 -3800
rect -936 -3864 -926 -3800
rect -794 -4322 -674 -3646
rect -103 -3877 -93 -3829
rect -329 -3977 -319 -3877
rect -267 -3929 -93 -3877
rect -41 -3929 -31 -3829
rect 42 -3929 52 -3829
rect 104 -3877 114 -3829
rect 104 -3929 252 -3877
rect -267 -3977 -257 -3929
rect 242 -3977 252 -3929
rect 304 -3977 314 -3877
rect 636 -3938 756 -3646
rect 1370 -3806 1380 -3729
rect 911 -3858 921 -3806
rect 1121 -3858 1380 -3806
rect 634 -3990 644 -3938
rect 744 -3990 756 -3938
rect -570 -4118 -560 -4062
rect -360 -4118 -350 -4062
rect 636 -4064 756 -3990
rect -103 -4187 -93 -4087
rect -41 -4135 -31 -4087
rect 636 -4116 646 -4064
rect 746 -4116 756 -4064
rect -41 -4187 252 -4135
rect 242 -4319 252 -4187
rect 304 -4319 314 -4135
rect -794 -4374 -784 -4322
rect -684 -4374 -674 -4322
rect -794 -4451 -674 -4374
rect 42 -4393 52 -4345
rect -795 -4503 -790 -4451
rect -685 -4503 -674 -4451
rect -329 -4493 -319 -4393
rect -267 -4445 52 -4393
rect 104 -4445 114 -4345
rect -267 -4493 -257 -4445
rect -1387 -4632 -1136 -4580
rect -936 -4632 -926 -4580
rect -1387 -6129 -1377 -4632
rect -794 -4713 -674 -4503
rect 335 -4638 345 -4574
rect 545 -4638 555 -4574
rect -797 -4765 -787 -4713
rect -687 -4765 -674 -4713
rect -794 -4838 -674 -4765
rect -794 -4890 -784 -4838
rect -684 -4890 -674 -4838
rect -1146 -5412 -1136 -5348
rect -936 -5412 -926 -5348
rect -794 -5870 -674 -4890
rect -103 -4909 -93 -4861
rect -329 -5034 -319 -4909
rect -267 -4961 -93 -4909
rect -41 -4961 -31 -4861
rect -267 -5034 -257 -4961
rect -570 -5150 -560 -5094
rect -360 -5150 -350 -5094
rect 636 -5096 756 -4116
rect 911 -4376 921 -4320
rect 1121 -4376 1131 -4320
rect 911 -4892 921 -4836
rect 1121 -4892 1131 -4836
rect 42 -5219 52 -5119
rect 104 -5167 114 -5119
rect 636 -5148 646 -5096
rect 746 -5148 756 -5096
rect 104 -5219 252 -5167
rect 242 -5267 252 -5219
rect 304 -5267 314 -5167
rect 636 -5230 756 -5148
rect 636 -5282 646 -5230
rect 746 -5282 756 -5230
rect 636 -5485 756 -5282
rect 1370 -5354 1380 -3858
rect 911 -5406 921 -5354
rect 1121 -5406 1380 -5354
rect 636 -5537 648 -5485
rect 748 -5537 758 -5485
rect -570 -5666 -560 -5610
rect -360 -5666 -350 -5610
rect 636 -5612 756 -5537
rect -103 -5735 -93 -5635
rect -41 -5683 -31 -5635
rect 636 -5664 646 -5612
rect 746 -5664 756 -5612
rect -41 -5735 252 -5683
rect 242 -5867 252 -5735
rect 304 -5867 314 -5683
rect -794 -5922 -784 -5870
rect -684 -5922 -674 -5870
rect -794 -6004 -674 -5922
rect 42 -5941 52 -5893
rect -795 -6056 -785 -6004
rect -685 -6056 -674 -6004
rect -329 -6041 -319 -5941
rect -267 -5993 52 -5941
rect 104 -5993 114 -5893
rect -267 -6041 -257 -5993
rect -1387 -6181 -1136 -6129
rect -936 -6181 -926 -6129
rect -1387 -7676 -1377 -6181
rect -794 -6256 -674 -6056
rect 335 -6186 345 -6122
rect 545 -6186 555 -6122
rect -794 -6308 -782 -6256
rect -682 -6308 -672 -6256
rect -794 -6386 -674 -6308
rect -794 -6438 -784 -6386
rect -684 -6438 -674 -6386
rect -1146 -6960 -1136 -6896
rect -936 -6960 -926 -6896
rect -794 -7418 -674 -6438
rect -103 -6457 -93 -6409
rect -329 -6583 -319 -6457
rect -267 -6509 -93 -6457
rect -41 -6509 -31 -6409
rect -267 -6583 -257 -6509
rect -570 -6698 -560 -6642
rect -360 -6698 -350 -6642
rect 636 -6644 756 -5664
rect 911 -5924 921 -5868
rect 1121 -5924 1131 -5868
rect 911 -6440 921 -6384
rect 1121 -6440 1131 -6384
rect 42 -6767 52 -6667
rect 104 -6715 114 -6667
rect 635 -6696 645 -6644
rect 745 -6696 756 -6644
rect 104 -6767 252 -6715
rect 242 -6815 252 -6767
rect 304 -6815 314 -6715
rect 636 -6781 756 -6696
rect 636 -6833 648 -6781
rect 748 -6833 758 -6781
rect 636 -7043 756 -6833
rect 1370 -6902 1380 -5406
rect 911 -6954 921 -6902
rect 1121 -6954 1380 -6902
rect 636 -7095 646 -7043
rect 746 -7095 756 -7043
rect -570 -7214 -560 -7158
rect -360 -7214 -350 -7158
rect 636 -7160 756 -7095
rect -103 -7283 -93 -7183
rect -41 -7231 -31 -7183
rect 636 -7212 646 -7160
rect 746 -7212 756 -7160
rect -41 -7283 252 -7231
rect 242 -7415 252 -7283
rect 304 -7415 314 -7231
rect -794 -7470 -784 -7418
rect -684 -7470 -674 -7418
rect -794 -7549 -674 -7470
rect 42 -7489 52 -7441
rect -794 -7601 -783 -7549
rect -683 -7601 -673 -7549
rect -329 -7589 -319 -7489
rect -267 -7541 52 -7489
rect 104 -7541 114 -7441
rect -267 -7589 -257 -7541
rect -1387 -7728 -1136 -7676
rect -936 -7728 -926 -7676
rect -1387 -9224 -1377 -7728
rect -794 -7811 -674 -7601
rect 335 -7734 345 -7670
rect 545 -7734 555 -7670
rect -795 -7863 -785 -7811
rect -685 -7863 -674 -7811
rect -794 -7934 -674 -7863
rect -794 -7986 -784 -7934
rect -684 -7986 -674 -7934
rect -1146 -8508 -1136 -8444
rect -936 -8508 -926 -8444
rect -794 -8966 -674 -7986
rect -103 -8005 -93 -7957
rect -329 -8131 -319 -8005
rect -267 -8057 -93 -8005
rect -41 -8057 -31 -7957
rect -267 -8131 -257 -8057
rect -329 -8137 -257 -8131
rect -570 -8246 -560 -8190
rect -360 -8246 -350 -8190
rect 636 -8192 756 -7212
rect 911 -7472 921 -7416
rect 1121 -7472 1131 -7416
rect 911 -7988 921 -7932
rect 1121 -7988 1131 -7932
rect 42 -8315 52 -8215
rect 104 -8263 114 -8215
rect 636 -8244 646 -8192
rect 746 -8244 756 -8192
rect 104 -8315 252 -8263
rect 242 -8363 252 -8315
rect 304 -8363 314 -8263
rect 636 -8329 756 -8244
rect 634 -8381 644 -8329
rect 744 -8381 756 -8329
rect 636 -8585 756 -8381
rect 1370 -8450 1380 -6954
rect 911 -8502 921 -8450
rect 1121 -8502 1380 -8450
rect 635 -8637 645 -8585
rect 745 -8637 756 -8585
rect -570 -8762 -560 -8706
rect -360 -8762 -350 -8706
rect 636 -8708 756 -8637
rect -103 -8831 -93 -8731
rect -41 -8779 -31 -8731
rect 636 -8760 646 -8708
rect 746 -8760 756 -8708
rect -41 -8831 252 -8779
rect -794 -9018 -784 -8966
rect -684 -9018 -674 -8966
rect 242 -8979 252 -8831
rect 304 -8979 314 -8779
rect -794 -9093 -674 -9018
rect 42 -9037 52 -8989
rect -794 -9145 -784 -9093
rect -684 -9145 -674 -9093
rect -329 -9137 -319 -9037
rect -267 -9089 52 -9037
rect 104 -9089 114 -8989
rect -267 -9137 -257 -9089
rect -1387 -9276 -1136 -9224
rect -936 -9276 -926 -9224
rect -1387 -10206 -1377 -9276
rect -794 -9358 -674 -9145
rect 335 -9282 345 -9218
rect 545 -9282 555 -9218
rect -794 -9410 -784 -9358
rect -684 -9410 -674 -9358
rect -794 -9482 -674 -9410
rect -794 -9534 -784 -9482
rect -684 -9534 -674 -9482
rect -103 -9553 -93 -9505
rect -329 -9653 -319 -9553
rect -267 -9605 -93 -9553
rect -41 -9605 -31 -9505
rect -267 -9653 -257 -9605
rect -570 -9794 -560 -9738
rect -360 -9794 -350 -9738
rect 636 -9740 756 -8760
rect 911 -9020 921 -8964
rect 1121 -9020 1131 -8964
rect 910 -9536 920 -9480
rect 1120 -9536 1130 -9480
rect 42 -9863 52 -9763
rect 104 -9811 114 -9763
rect 636 -9792 646 -9740
rect 746 -9792 756 -9740
rect 104 -9863 252 -9811
rect 242 -9911 252 -9863
rect 304 -9911 314 -9811
rect 636 -9863 756 -9792
rect 636 -9915 648 -9863
rect 748 -9915 758 -9863
rect 636 -9939 756 -9915
rect -1146 -10056 -1136 -9992
rect -936 -10056 -926 -9992
rect 1370 -9998 1380 -8502
rect 911 -10050 921 -9998
rect 1121 -10050 1380 -9998
rect 1370 -10070 1380 -10050
rect 1492 -9045 1502 -3729
rect 2112 -8325 2122 -2918
rect 2313 -8325 2323 -2918
rect 2962 -2936 3062 -2807
rect 2962 -2988 3269 -2936
rect 3392 -2988 3402 -2936
rect 2962 -3001 3062 -2988
rect 2472 -3053 2482 -3001
rect 2542 -3053 2598 -3001
rect 2658 -3053 3062 -3001
rect 2472 -3517 2552 -3053
rect 2472 -3569 2482 -3517
rect 2542 -3569 2552 -3517
rect 2472 -4033 2552 -3569
rect 2588 -3311 2598 -3259
rect 2658 -3311 2668 -3259
rect 2588 -3517 2668 -3311
rect 3700 -3394 3710 -2888
rect 3312 -3446 3322 -3394
rect 3445 -3446 3710 -3394
rect 2588 -3569 3269 -3517
rect 3392 -3569 3401 -3517
rect 2588 -3775 2668 -3569
rect 2588 -3827 2598 -3775
rect 2658 -3827 2668 -3775
rect 3700 -3975 3710 -3446
rect 3311 -4027 3321 -3975
rect 3445 -4027 3710 -3975
rect 2472 -4085 2482 -4033
rect 2542 -4085 2552 -4033
rect 3700 -4242 3710 -4027
rect 3861 -4242 3871 -2888
rect 2472 -4343 2482 -4291
rect 2542 -4343 2552 -4291
rect 2472 -4807 2552 -4343
rect 2472 -4859 2482 -4807
rect 2542 -4859 2552 -4807
rect 2472 -5323 2552 -4859
rect 2588 -4601 2598 -4549
rect 2658 -4601 2668 -4549
rect 2588 -4807 2668 -4601
rect 2588 -4859 3269 -4807
rect 3382 -4859 3392 -4807
rect 2588 -5065 2668 -4859
rect 2588 -5117 2598 -5065
rect 2658 -5117 2668 -5065
rect 3706 -5265 3716 -4242
rect 3312 -5317 3322 -5265
rect 3445 -5317 3716 -5265
rect 2472 -5375 2482 -5323
rect 2542 -5375 2552 -5323
rect 2472 -5633 2482 -5581
rect 2542 -5633 2552 -5581
rect 2472 -6097 2552 -5633
rect 2472 -6149 2482 -6097
rect 2542 -6149 2552 -6097
rect 2472 -6607 2552 -6149
rect 2588 -5891 2598 -5839
rect 2658 -5891 2668 -5839
rect 2588 -6097 2668 -5891
rect 2588 -6149 3269 -6097
rect 3382 -6149 3392 -6097
rect 2588 -6355 2668 -6149
rect 2588 -6407 2598 -6355
rect 2658 -6407 2668 -6355
rect 3706 -6555 3716 -5317
rect 3312 -6607 3322 -6555
rect 3445 -6607 3716 -6555
rect 2472 -6671 2482 -6607
rect 2546 -6671 2556 -6607
rect 2472 -6923 2482 -6871
rect 2542 -6923 2552 -6871
rect 2472 -7387 2552 -6923
rect 2472 -7439 2482 -7387
rect 2542 -7439 2552 -7387
rect 2472 -7903 2552 -7439
rect 2588 -7181 2598 -7129
rect 2658 -7181 2668 -7129
rect 2588 -7387 2668 -7181
rect 2588 -7439 3269 -7387
rect 3382 -7439 3392 -7387
rect 2588 -7645 2668 -7439
rect 2588 -7697 2598 -7645
rect 2658 -7697 2668 -7645
rect 3706 -7845 3716 -6607
rect 3312 -7897 3322 -7845
rect 3445 -7895 3716 -7845
rect 3855 -7254 3865 -4242
rect 6757 -6606 6836 111
rect 7148 108 7183 115
rect 7148 105 11593 108
rect 7183 98 11593 105
rect 8506 -25 10634 -15
rect 8564 -138 10634 -128
rect 9080 -293 9132 -292
rect 9996 -293 10048 -292
rect 9080 -302 10928 -293
rect 9132 -393 9996 -302
rect 9080 -472 9132 -462
rect 10048 -393 10928 -302
rect 9518 -473 9612 -463
rect 9996 -472 10048 -462
rect 9518 -620 9612 -610
rect 8506 -676 8564 -666
rect 8599 -731 8693 -721
rect 8599 -878 8693 -868
rect 10434 -731 10528 -721
rect 10434 -878 10528 -868
rect 8861 -919 9061 -909
rect 8861 -981 9061 -971
rect 9319 -919 9519 -909
rect 9319 -981 9519 -971
rect 9777 -919 9977 -909
rect 9777 -981 9977 -971
rect 10235 -919 10435 -909
rect 10235 -981 10435 -971
rect 7122 -1043 7205 -1033
rect 7122 -1153 7205 -1143
rect 8961 -1043 9061 -981
rect 8961 -1153 9061 -1143
rect 9151 -1043 9251 -1033
rect 7112 -1229 7225 -1219
rect 7112 -1339 7225 -1329
rect 8693 -1229 8793 -1219
rect 8693 -1406 8793 -1329
rect 9151 -1406 9251 -1143
rect 9419 -1229 9519 -981
rect 9419 -1339 9519 -1329
rect 9609 -1043 9709 -1033
rect 9609 -1406 9709 -1143
rect 9877 -1229 9977 -981
rect 10335 -1043 10435 -981
rect 10335 -1153 10435 -1143
rect 9877 -1339 9977 -1329
rect 10067 -1229 10167 -1219
rect 10067 -1406 10167 -1329
rect 8693 -1416 8893 -1406
rect 8693 -1478 8893 -1468
rect 9151 -1416 9351 -1406
rect 9151 -1478 9351 -1468
rect 9609 -1416 9809 -1406
rect 9609 -1478 9809 -1468
rect 10067 -1416 10267 -1406
rect 10067 -1478 10267 -1468
rect 8600 -1520 8694 -1510
rect 8600 -1667 8694 -1657
rect 10432 -1520 10526 -1510
rect 10432 -1667 10526 -1657
rect 8497 -1702 8571 -1692
rect 7733 -1785 8045 -1775
rect 8045 -2003 8497 -1785
rect 7733 -2013 8045 -2003
rect 8452 -2333 8497 -2323
rect 9517 -1731 9611 -1721
rect 9517 -1878 9611 -1868
rect 9080 -1925 9132 -1915
rect 9996 -1925 10048 -1915
rect 9132 -2085 9996 -1992
rect 10828 -1992 10928 -393
rect 11697 -420 12178 -410
rect 11697 -552 11770 -420
rect 11822 -552 12126 -420
rect 11770 -630 11822 -620
rect 12126 -630 12178 -620
rect 11593 -1061 11697 -1051
rect 11898 -716 11950 -706
rect 11898 -1302 11950 -916
rect 11898 -1391 11950 -1381
rect 12254 -716 12306 -706
rect 12254 -1136 12306 -916
rect 12254 -1316 14187 -1136
rect 12254 -1425 12306 -1316
rect 12254 -1506 12306 -1496
rect 11810 -1530 11862 -1520
rect 11810 -1875 11862 -1601
rect 12166 -1530 12218 -1520
rect 12166 -1875 12218 -1601
rect 10048 -2085 10928 -1992
rect 9080 -2092 10928 -2085
rect 10997 -1885 12375 -1875
rect 9080 -2095 9132 -2092
rect 9996 -2095 10127 -2092
rect 8571 -2330 8679 -2323
rect 8571 -2333 9795 -2330
rect 8679 -2340 9795 -2333
rect 8410 -3760 8452 -3486
rect 8790 -2520 9795 -2510
rect 10005 -2609 10127 -2095
rect 10997 -2167 12375 -2157
rect 11087 -2367 11228 -2357
rect 11228 -2377 11495 -2367
rect 12537 -2368 12609 -1316
rect 11228 -2429 11293 -2377
rect 11087 -2439 11228 -2429
rect 11293 -2439 11495 -2429
rect 12127 -2378 12609 -2368
rect 12329 -2430 12609 -2378
rect 12127 -2440 12609 -2430
rect 10341 -2468 10552 -2458
rect 9719 -2619 10128 -2609
rect 9719 -2694 10128 -2684
rect 8957 -2712 9013 -2702
rect 8957 -2862 9013 -2852
rect 8790 -2978 9552 -2968
rect 8790 -3042 9052 -2978
rect 8790 -3052 9552 -3042
rect 10005 -3325 10127 -2694
rect 9719 -3335 10128 -3325
rect 9719 -3410 10128 -3400
rect 8790 -3519 10341 -3509
rect 8679 -3760 10341 -3758
rect 8410 -3768 10341 -3760
rect 8410 -3770 8679 -3768
rect 8410 -3771 8570 -3770
rect 10341 -3779 10552 -3769
rect 6757 -6682 6836 -6672
rect 4485 -7254 4907 -7244
rect 3855 -7642 4485 -7254
rect 3855 -7895 3865 -7642
rect 4485 -7652 4907 -7642
rect 3445 -7897 3865 -7895
rect 2472 -7955 2482 -7903
rect 2542 -7955 2552 -7903
rect 2112 -8418 2323 -8325
rect 2472 -8213 2482 -8161
rect 2542 -8213 2552 -8161
rect 2472 -8579 2552 -8213
rect 3706 -8356 3865 -7897
rect 3706 -8357 3815 -8356
rect 3259 -8533 3269 -8469
rect 3409 -8533 3419 -8469
rect 1750 -8659 1760 -8579
rect 1833 -8659 2552 -8579
rect 3592 -8733 3602 -8357
rect 3295 -8785 3305 -8733
rect 3445 -8785 3602 -8733
rect 1492 -9069 2893 -9045
rect 3259 -9049 3269 -8985
rect 3409 -9049 3419 -8985
rect 1492 -9177 1720 -9069
rect 2763 -9177 2893 -9069
rect 1492 -9199 2893 -9177
rect 1492 -9551 1502 -9199
rect 2703 -9302 2893 -9199
rect 1956 -9444 1966 -9370
rect 2566 -9444 2576 -9370
rect 1492 -10070 1541 -9551
rect 1370 -10078 1541 -10070
rect 1637 -10078 1647 -9551
rect 2703 -10078 2730 -9302
rect 1370 -10083 1647 -10078
rect 1370 -10206 1424 -10083
rect -1387 -10260 -1305 -10206
rect -1153 -10260 -315 -10206
rect -167 -10260 1424 -10206
rect 2141 -10104 2730 -10078
rect 2141 -10224 2153 -10104
rect 2632 -10127 2730 -10104
rect 2878 -10127 2893 -9302
rect 3139 -9636 3149 -9277
rect 3214 -9636 3224 -9277
rect 3592 -9343 3602 -8785
rect 3737 -9343 3815 -8357
rect 3594 -9658 3604 -9343
rect 3259 -9710 3269 -9658
rect 3345 -9710 3604 -9658
rect 3139 -10090 3149 -9731
rect 3214 -10090 3224 -9731
rect 3594 -9918 3604 -9710
rect 3575 -9970 3604 -9918
rect 2632 -10224 2893 -10127
rect 2141 -10239 2893 -10224
rect -1387 -10263 -1377 -10260
rect -1571 -10375 -1377 -10263
rect 3594 -10336 3604 -9970
rect 3736 -10335 3815 -9343
rect 3963 -10335 3973 -8356
rect 3736 -10336 3973 -10335
rect 3660 -10337 3973 -10336
rect 3809 -10407 3973 -10337
<< via2 >>
rect -1749 7491 730 7598
rect -10065 1687 -9489 1697
rect -10065 1632 -9489 1687
rect -9450 640 -9447 1438
rect -9447 640 -9395 1438
rect -9395 640 -9392 1438
rect -615 5392 -551 6392
rect -1492 4155 -1428 5155
rect 261 4155 325 5155
rect -6292 2358 -6236 2371
rect -6292 2039 -6288 2358
rect -6288 2039 -6236 2358
rect -6292 2029 -6236 2039
rect -6293 1277 -6235 1287
rect -6293 958 -6289 1277
rect -6289 958 -6237 1277
rect -6237 958 -6235 1277
rect -6293 948 -6235 958
rect -10599 -266 -10501 134
rect -8677 89 -8197 92
rect -8677 37 -8197 89
rect -8677 34 -8197 37
rect -6219 90 -5739 94
rect -6219 38 -5739 90
rect -6219 36 -5739 38
rect -1491 2154 -1427 3154
rect 261 2154 325 3154
rect -615 994 -551 1994
rect 1715 3760 1725 3860
rect 1725 3760 2007 3860
rect 7431 1669 7495 1869
rect 9547 1945 9611 2145
rect 11663 1669 11727 1869
rect 13414 2399 13712 2786
rect 7431 783 7495 983
rect 9547 507 9611 707
rect 11663 783 11727 983
rect -1481 -972 -1417 -872
rect 6271 -972 6335 -872
rect 2395 -1148 2459 -1048
rect 2395 -1382 2459 -1282
rect -1481 -1558 -1417 -1458
rect 6271 -1558 6335 -1458
rect 6245 -2003 6429 -1786
rect 2962 -2494 3062 -2314
rect 2962 -2807 3062 -2707
rect -1136 -3864 -936 -3800
rect -560 -4118 -360 -4062
rect 345 -4638 545 -4574
rect -1136 -5412 -936 -5348
rect -560 -5150 -360 -5094
rect 921 -4376 1121 -4320
rect 921 -4892 1121 -4836
rect -560 -5666 -360 -5610
rect 345 -6186 545 -6122
rect -1136 -6960 -936 -6896
rect -560 -6698 -360 -6642
rect 921 -5924 1121 -5868
rect 921 -6440 1121 -6384
rect -560 -7214 -360 -7158
rect 345 -7734 545 -7670
rect -1136 -8508 -936 -8444
rect -560 -8246 -360 -8190
rect 921 -7472 1121 -7416
rect 921 -7988 1121 -7932
rect -560 -8762 -360 -8706
rect 345 -9282 545 -9218
rect -560 -9794 -360 -9738
rect 921 -9020 1121 -8964
rect 920 -9536 1120 -9480
rect -1136 -10056 -936 -9992
rect 2482 -6613 2546 -6607
rect 2482 -6665 2542 -6613
rect 2542 -6665 2546 -6613
rect 2482 -6671 2546 -6665
rect 9518 -610 9612 -473
rect 8599 -868 8693 -731
rect 10434 -868 10528 -731
rect 7122 -1143 7205 -1043
rect 7112 -1329 7225 -1229
rect 8600 -1657 8694 -1520
rect 10432 -1657 10526 -1520
rect 7733 -2003 8045 -1785
rect 9517 -1868 9611 -1731
rect 11087 -2429 11228 -2367
rect 8957 -2852 9013 -2712
rect 6757 -6672 6836 -6606
rect 4485 -7642 4907 -7254
rect 3269 -8533 3409 -8469
rect 1760 -8659 1833 -8579
rect 3269 -9049 3409 -8985
rect 1966 -9444 2566 -9370
rect 3149 -9636 3214 -9277
rect 3149 -10090 3214 -9731
<< metal3 >>
rect -1759 7598 740 7603
rect -1759 7491 -1749 7598
rect 730 7491 740 7598
rect -1759 7486 740 7491
rect -625 6392 -541 6397
rect -625 5392 -615 6392
rect -551 5478 -541 6392
rect 2950 5893 5030 5913
rect 2950 5829 2978 5893
rect 5002 5829 5030 5893
rect -551 5392 567 5478
rect -625 5387 567 5392
rect -611 5378 567 5387
rect -1502 5155 -1418 5160
rect -1502 4155 -1492 5155
rect -1428 4155 -1418 5155
rect -1502 4150 -1418 4155
rect 251 5155 335 5160
rect 251 4155 261 5155
rect 325 4155 335 5155
rect 251 4150 335 4155
rect 467 3162 567 5378
rect 2950 4562 5030 5829
rect 2950 4382 13000 4562
rect 2950 3865 5030 4382
rect 1705 3860 5030 3865
rect 1705 3760 1715 3860
rect 2007 3760 5030 3860
rect 1705 3755 5030 3760
rect 2950 3541 5030 3755
rect 467 3159 658 3162
rect -1501 3154 658 3159
rect -6303 2371 -6225 2376
rect -6303 2029 -6292 2371
rect -6236 2029 -6225 2371
rect -1501 2154 -1491 3154
rect -1427 3059 261 3154
rect -1427 2154 -1417 3059
rect -1501 2149 -1417 2154
rect 251 2154 261 3059
rect 325 3059 658 3154
rect 325 2154 335 3059
rect 251 2149 335 2154
rect -6303 1702 -6225 2029
rect -10075 1697 -6225 1702
rect -10075 1632 -10065 1697
rect -9489 1632 -6225 1697
rect -10075 1627 -6225 1632
rect -9460 1438 -9280 1443
rect -9460 640 -9450 1438
rect -9392 640 -9280 1438
rect -6303 1287 -6225 1627
rect -6303 948 -6293 1287
rect -6235 948 -6225 1287
rect -625 1994 -541 1999
rect -625 994 -615 1994
rect -551 994 -541 1994
rect -625 989 -541 994
rect -6303 943 -6225 948
rect -10609 134 -10491 139
rect -10609 -266 -10599 134
rect -10501 -266 -10491 134
rect -10609 -271 -10491 -266
rect -9460 -326 -9280 640
rect -8687 92 -8187 97
rect -8687 34 -8677 92
rect -8197 34 -8187 92
rect -8687 29 -8187 34
rect -6229 94 -5729 99
rect -6229 36 -6219 94
rect -5739 36 -5729 94
rect -6229 31 -5729 36
rect -9470 -430 -9460 -326
rect -9280 -430 -9270 -326
rect -9460 -525 -9280 -430
rect -8687 -991 -8507 29
rect -6229 -958 -6049 31
rect -1498 -872 -1400 -867
rect -1498 -972 -1481 -872
rect -1417 -972 -1400 -872
rect -1498 -977 -1400 -972
rect 548 -1043 658 3059
rect 9537 2145 9621 2150
rect 9537 1945 9547 2145
rect 9611 1945 9621 2145
rect 9537 1940 9621 1945
rect 7421 1869 7505 1874
rect 7421 1669 7431 1869
rect 7495 1764 7505 1869
rect 11653 1869 11737 1874
rect 11653 1764 11663 1869
rect 7495 1669 11663 1764
rect 11727 1764 11737 1869
rect 11727 1669 12177 1764
rect 7421 1664 12177 1669
rect 7421 983 7505 988
rect 7421 783 7431 983
rect 7495 783 7505 983
rect 7421 778 7505 783
rect 11653 983 11737 988
rect 11653 783 11663 983
rect 11727 783 11737 983
rect 11653 778 11737 783
rect 9537 707 9621 712
rect 9537 507 9547 707
rect 9611 602 9621 707
rect 12077 602 12177 1664
rect 9611 507 12177 602
rect 9537 502 12177 507
rect 9508 -473 9622 -468
rect 9508 -610 9518 -473
rect 9612 -610 9622 -473
rect 9508 -615 9622 -610
rect 10707 -726 10854 502
rect 8589 -731 10854 -726
rect 6233 -872 6361 -867
rect 6233 -972 6271 -872
rect 6335 -972 6361 -872
rect 8589 -868 8599 -731
rect 8693 -868 10434 -731
rect 10528 -868 10854 -731
rect 8589 -873 10854 -868
rect 6233 -977 6361 -972
rect 7112 -1043 7215 -1038
rect 548 -1048 6731 -1043
rect 548 -1148 2395 -1048
rect 2459 -1148 6731 -1048
rect 7081 -1143 7122 -1043
rect 7205 -1143 7215 -1043
rect 7112 -1148 7215 -1143
rect 548 -1153 6731 -1148
rect 6621 -1229 6731 -1153
rect 7102 -1229 7235 -1224
rect 2369 -1282 2484 -1277
rect 2369 -1382 2395 -1282
rect 2459 -1382 2484 -1282
rect 2369 -1387 2484 -1382
rect 6621 -1329 7112 -1229
rect 7225 -1329 7235 -1229
rect 6621 -1453 6731 -1329
rect 7102 -1334 7235 -1329
rect -1491 -1458 6731 -1453
rect -1491 -1558 -1481 -1458
rect -1417 -1558 6271 -1458
rect 6335 -1558 6731 -1458
rect -1491 -1563 6731 -1558
rect 8590 -1520 8704 -1515
rect 8590 -1657 8600 -1520
rect 8694 -1657 8704 -1520
rect 8590 -1662 8704 -1657
rect 10422 -1520 10536 -1515
rect 10422 -1657 10432 -1520
rect 10526 -1657 10536 -1520
rect 10422 -1662 10536 -1657
rect 9507 -1731 9621 -1726
rect 10707 -1731 10854 -873
rect 6235 -1786 6439 -1781
rect 6235 -2003 6245 -1786
rect 6429 -2003 6439 -1786
rect 6235 -2008 6439 -2003
rect 7723 -1785 8055 -1780
rect 7723 -2003 7733 -1785
rect 8045 -2003 8055 -1785
rect 9507 -1868 9517 -1731
rect 9611 -1868 10854 -1731
rect 9507 -1873 10854 -1868
rect 7723 -2008 8055 -2003
rect 2952 -2314 3072 -2309
rect 2952 -2494 2962 -2314
rect 3062 -2494 3072 -2314
rect 11077 -2364 11238 -2362
rect 11077 -2432 11087 -2364
rect 11228 -2432 11238 -2364
rect 11077 -2434 11238 -2432
rect 2952 -2499 3072 -2494
rect 2952 -2707 3072 -2702
rect 2952 -2807 2962 -2707
rect 3062 -2712 9023 -2707
rect 3062 -2807 8957 -2712
rect 2952 -2812 3072 -2807
rect 8947 -2852 8957 -2807
rect 9013 -2852 9023 -2712
rect 8947 -2857 9023 -2852
rect 12820 -2953 13000 4382
rect 13404 2786 13722 2791
rect 13404 2399 13414 2786
rect 13712 2399 13722 2786
rect 13404 2394 13722 2399
rect 10789 -2981 14561 -2953
rect -1141 -3800 -931 -3790
rect -1141 -3864 -1136 -3800
rect -936 -3864 -931 -3800
rect -1141 -3874 -931 -3864
rect 10789 -3926 14477 -2981
rect 10567 -4033 14477 -3926
rect -565 -4062 -355 -4052
rect -565 -4118 -560 -4062
rect -360 -4118 -355 -4062
rect -565 -4128 -355 -4118
rect -431 -4192 -355 -4128
rect -431 -5084 -357 -4192
rect 916 -4320 1126 -4310
rect 916 -4376 921 -4320
rect 1121 -4376 1126 -4320
rect 916 -4386 1126 -4376
rect 340 -4574 550 -4564
rect 340 -4638 345 -4574
rect 545 -4638 550 -4574
rect 340 -4648 550 -4638
rect 1050 -4826 1126 -4386
rect 916 -4836 1126 -4826
rect 916 -4892 921 -4836
rect 1121 -4892 1126 -4836
rect 916 -4902 1126 -4892
rect -565 -5094 -355 -5084
rect -565 -5150 -560 -5094
rect -360 -5150 -355 -5094
rect -565 -5160 -355 -5150
rect -1141 -5348 -931 -5338
rect -1141 -5412 -1136 -5348
rect -936 -5412 -931 -5348
rect -1141 -5422 -931 -5412
rect -431 -5600 -357 -5160
rect -565 -5610 -355 -5600
rect -565 -5666 -560 -5610
rect -360 -5666 -355 -5610
rect -565 -5676 -355 -5666
rect -431 -6632 -357 -5676
rect 1050 -5858 1126 -4902
rect 916 -5868 1126 -5858
rect 916 -5924 921 -5868
rect 1121 -5924 1126 -5868
rect 916 -5934 1126 -5924
rect 340 -6122 550 -6112
rect 340 -6186 345 -6122
rect 545 -6186 550 -6122
rect 340 -6196 550 -6186
rect 1050 -6374 1126 -5934
rect 916 -6384 1126 -6374
rect 916 -6440 921 -6384
rect 1121 -6440 1126 -6384
rect 10789 -6405 14477 -4033
rect 14541 -6405 14561 -2981
rect 10789 -6433 14561 -6405
rect 916 -6450 1126 -6440
rect -565 -6642 -355 -6632
rect -565 -6698 -560 -6642
rect -360 -6698 -355 -6642
rect -565 -6708 -355 -6698
rect -1141 -6896 -931 -6886
rect -1141 -6960 -1136 -6896
rect -936 -6960 -931 -6896
rect -1141 -6970 -931 -6960
rect -431 -7148 -357 -6708
rect -565 -7158 -355 -7148
rect -565 -7214 -560 -7158
rect -360 -7214 -355 -7158
rect -565 -7224 -355 -7214
rect -431 -8180 -357 -7224
rect 1050 -7406 1126 -6450
rect 2477 -6607 2594 -6597
rect 2477 -6671 2482 -6607
rect 2546 -6671 2594 -6607
rect 2477 -6681 2594 -6671
rect 6730 -6606 6853 -6599
rect 6730 -6672 6757 -6606
rect 6836 -6672 6853 -6606
rect 6730 -6683 6853 -6672
rect 916 -7416 1126 -7406
rect 916 -7472 921 -7416
rect 1121 -7472 1126 -7416
rect 916 -7482 1126 -7472
rect 340 -7670 550 -7660
rect 340 -7734 345 -7670
rect 545 -7734 550 -7670
rect 340 -7744 550 -7734
rect 1050 -7922 1126 -7482
rect 4475 -7254 4917 -7249
rect 4475 -7642 4485 -7254
rect 4907 -7642 4917 -7254
rect 4475 -7647 4917 -7642
rect 916 -7932 1126 -7922
rect 916 -7988 921 -7932
rect 1121 -7988 1126 -7932
rect 916 -7998 1126 -7988
rect -565 -8190 -355 -8180
rect -565 -8246 -560 -8190
rect -360 -8246 -355 -8190
rect -565 -8256 -355 -8246
rect -1141 -8444 -931 -8434
rect -1141 -8508 -1136 -8444
rect -936 -8508 -931 -8444
rect -1141 -8518 -931 -8508
rect -431 -8696 -357 -8256
rect -565 -8706 -355 -8696
rect -565 -8762 -560 -8706
rect -360 -8762 -355 -8706
rect -565 -8772 -355 -8762
rect -431 -9728 -357 -8772
rect 1050 -8878 1126 -7998
rect 3264 -8469 3414 -8459
rect 3264 -8533 3269 -8469
rect 3409 -8533 3414 -8469
rect 3264 -8543 3414 -8533
rect 1755 -8579 1838 -8569
rect 1755 -8659 1760 -8579
rect 1833 -8659 1838 -8579
rect 1755 -8669 1838 -8659
rect 1760 -8878 1833 -8669
rect 1050 -8954 1833 -8878
rect 916 -8964 1126 -8954
rect 916 -9020 921 -8964
rect 1121 -9020 1126 -8964
rect 916 -9030 1126 -9020
rect 340 -9218 550 -9208
rect 340 -9282 345 -9218
rect 545 -9282 550 -9218
rect 340 -9292 550 -9282
rect 1050 -9470 1126 -9030
rect 3264 -8985 3414 -8975
rect 3264 -9049 3269 -8985
rect 3409 -9049 3414 -8985
rect 3264 -9059 3414 -9049
rect 3144 -9277 3219 -9267
rect 1961 -9370 2571 -9360
rect 1961 -9444 1966 -9370
rect 2566 -9444 2571 -9370
rect 1961 -9454 2571 -9444
rect 915 -9480 1126 -9470
rect 915 -9536 920 -9480
rect 1120 -9536 1126 -9480
rect 915 -9546 1126 -9536
rect -565 -9738 -355 -9728
rect -565 -9794 -560 -9738
rect -360 -9794 -355 -9738
rect -565 -9804 -355 -9794
rect -1141 -9992 -931 -9982
rect -1141 -10056 -1136 -9992
rect -936 -10056 -931 -9992
rect -1141 -10066 -931 -10056
rect -431 -10120 -357 -9804
rect 1050 -10120 1126 -9546
rect 3144 -9636 3149 -9277
rect 3214 -9636 3219 -9277
rect 3144 -9646 3219 -9636
rect 3144 -9731 3219 -9721
rect 3144 -10090 3149 -9731
rect 3214 -10090 3219 -9731
rect 3144 -10100 3219 -10090
rect -431 -10194 1126 -10120
<< via3 >>
rect -1749 7491 730 7598
rect 2978 5829 5002 5893
rect -1492 4155 -1428 5155
rect 261 4155 325 5155
rect -615 994 -551 1994
rect -10599 -266 -10501 134
rect -9460 -430 -9280 -326
rect -1481 -972 -1417 -872
rect 9547 1945 9611 2145
rect 7431 783 7495 983
rect 11663 783 11727 983
rect 9518 -610 9612 -473
rect 6271 -972 6335 -872
rect 7122 -1143 7205 -1043
rect 2395 -1382 2459 -1282
rect 7112 -1329 7225 -1229
rect 8600 -1657 8694 -1520
rect 10432 -1657 10526 -1520
rect 6245 -2003 6429 -1786
rect 7733 -2003 8045 -1785
rect 2962 -2494 3062 -2314
rect 11087 -2367 11228 -2364
rect 11087 -2429 11228 -2367
rect 11087 -2432 11228 -2429
rect 13414 2399 13712 2786
rect -1136 -3864 -936 -3800
rect 345 -4638 545 -4574
rect -1136 -5412 -936 -5348
rect 345 -6186 545 -6122
rect 14477 -6405 14541 -2981
rect -1136 -6960 -936 -6896
rect 2482 -6671 2546 -6607
rect 6757 -6672 6836 -6606
rect 345 -7734 545 -7670
rect 4485 -7642 4907 -7254
rect -1136 -8508 -936 -8444
rect 3269 -8533 3409 -8469
rect 345 -9282 545 -9218
rect 3269 -9049 3409 -8985
rect 1966 -9444 2566 -9370
rect -1136 -10056 -936 -9992
rect 3149 -9636 3214 -9277
rect 3149 -10090 3214 -9731
<< mimcap >>
rect 2990 5541 4990 5581
rect 2990 3621 3030 5541
rect 4950 3621 4990 5541
rect 2990 3581 4990 3621
rect 10829 -3033 14229 -2993
rect 10829 -6353 10869 -3033
rect 14189 -6353 14229 -3033
rect 10829 -6393 14229 -6353
<< mimcapcontact >>
rect 3030 3621 4950 5541
rect 10869 -6353 14189 -3033
<< metal4 >>
rect -1903 7598 897 7813
rect -1903 7491 -1749 7598
rect 730 7491 897 7598
rect -1903 7413 897 7491
rect 2962 5893 5018 5909
rect 2962 5829 2978 5893
rect 5002 5829 5018 5893
rect 2962 5813 5018 5829
rect 3029 5541 4951 5542
rect -1493 5155 -1427 5156
rect -1493 4155 -1492 5155
rect -1428 4254 -1427 5155
rect 260 5155 326 5156
rect 260 4254 261 5155
rect -1428 4155 261 4254
rect 325 4254 326 5155
rect 325 4155 961 4254
rect -1493 4154 961 4155
rect -616 1994 -550 1995
rect -616 994 -615 1994
rect -551 1960 -550 1994
rect 861 1960 961 4154
rect 3029 3621 3030 5541
rect 4950 3725 4951 5541
rect 4950 3659 6353 3725
rect 4950 3621 4951 3659
rect 3029 3620 4951 3621
rect -551 1860 961 1960
rect 6287 1946 6353 3659
rect 13413 2786 13713 2787
rect 13151 2399 13414 2786
rect 13712 2399 15660 2786
rect 13413 2398 13713 2399
rect -551 994 -550 1860
rect -616 993 -550 994
rect -10600 134 -10500 135
rect -10693 -266 -10599 134
rect -10501 -266 -10425 134
rect -10600 -267 -10500 -266
rect -9461 -326 -9279 -325
rect -9461 -430 -9460 -326
rect -9280 -430 -9279 -326
rect -9461 -431 -9279 -430
rect -9460 -548 -9280 -431
rect -9460 -728 -3326 -548
rect -3506 -2314 -3326 -728
rect 861 -871 961 1860
rect 6286 1868 6353 1946
rect 6978 2145 9612 2146
rect 6978 2046 9547 2145
rect 6286 -871 6352 1868
rect 6978 984 7078 2046
rect 9546 1945 9547 2046
rect 9611 1945 9612 2145
rect 9546 1944 9612 1945
rect 6978 983 11728 984
rect 6978 884 7431 983
rect 7430 783 7431 884
rect 7495 884 11663 983
rect 7495 783 7496 884
rect 7430 782 7496 783
rect 8323 -472 8462 884
rect 11662 783 11663 884
rect 11727 783 11728 983
rect 11662 782 11728 783
rect 8323 -473 9635 -472
rect 8323 -610 9518 -473
rect 9612 -610 9635 -473
rect 8323 -611 9635 -610
rect -1482 -872 6999 -871
rect -1482 -972 -1481 -872
rect -1417 -972 6271 -872
rect 6335 -972 6999 -872
rect -1482 -973 6999 -972
rect 6897 -1043 6999 -973
rect 7121 -1043 7206 -1042
rect 6897 -1143 7122 -1043
rect 7205 -1143 7206 -1043
rect 6897 -1281 6999 -1143
rect 7121 -1144 7206 -1143
rect 7111 -1229 7226 -1228
rect 2394 -1282 6999 -1281
rect 2394 -1382 2395 -1282
rect 2459 -1382 6999 -1282
rect 7087 -1329 7112 -1229
rect 7225 -1329 7226 -1229
rect 7111 -1330 7226 -1329
rect 2394 -1383 6999 -1382
rect 8323 -1519 8462 -611
rect 8323 -1520 10527 -1519
rect 8323 -1657 8600 -1520
rect 8694 -1657 10432 -1520
rect 10526 -1657 10527 -1520
rect 8323 -1658 10527 -1657
rect 7732 -1785 8046 -1784
rect 6244 -1786 7733 -1785
rect 6059 -2003 6245 -1786
rect 6429 -2003 7733 -1786
rect 8045 -2003 8517 -1785
rect 6244 -2004 6430 -2003
rect 7732 -2004 8046 -2003
rect 2961 -2314 3063 -2313
rect -3506 -2494 2962 -2314
rect 3062 -2494 3073 -2314
rect 11078 -2364 11229 -2363
rect 11078 -2432 11087 -2364
rect 11228 -2367 11229 -2364
rect 11228 -2429 11297 -2367
rect 11228 -2432 11229 -2429
rect 11078 -2433 11229 -2432
rect 2961 -2495 3063 -2494
rect 11078 -3032 11189 -2433
rect 14461 -2981 14557 -2965
rect 10868 -3033 14190 -3032
rect -1137 -3800 -935 -3799
rect -1137 -3864 -1136 -3800
rect -936 -3864 -935 -3800
rect -1137 -3865 -935 -3864
rect -1137 -5347 -1061 -3865
rect 344 -4574 546 -4573
rect 344 -4638 345 -4574
rect 545 -4638 546 -4574
rect 344 -4639 546 -4638
rect -1137 -5348 -935 -5347
rect -1137 -5412 -1136 -5348
rect -936 -5412 -935 -5348
rect -1137 -5413 -935 -5412
rect -1137 -6895 -1061 -5413
rect 344 -6121 420 -4639
rect 344 -6122 546 -6121
rect 344 -6186 345 -6122
rect 545 -6186 546 -6122
rect 344 -6187 546 -6186
rect -1137 -6896 -935 -6895
rect -1137 -6960 -1136 -6896
rect -936 -6960 -935 -6896
rect -1137 -6961 -935 -6960
rect -1137 -8443 -1061 -6961
rect 344 -7669 420 -6187
rect 10868 -6353 10869 -3033
rect 14189 -6353 14190 -3033
rect 10868 -6354 14190 -6353
rect 14461 -6405 14477 -2981
rect 14541 -6405 14557 -2981
rect 14461 -6421 14557 -6405
rect 6756 -6606 6837 -6605
rect 2481 -6607 6757 -6606
rect 2481 -6671 2482 -6607
rect 2546 -6671 6757 -6607
rect 2481 -6672 6757 -6671
rect 6836 -6672 6837 -6606
rect 6756 -6673 6837 -6672
rect 4484 -7254 4908 -7253
rect 15273 -7254 15660 2399
rect 4484 -7642 4485 -7254
rect 4907 -7641 15660 -7254
rect 4907 -7642 4908 -7641
rect 4484 -7643 4908 -7642
rect 344 -7670 546 -7669
rect 344 -7734 345 -7670
rect 545 -7734 546 -7670
rect 344 -7735 546 -7734
rect -1137 -8444 -935 -8443
rect -1137 -8508 -1136 -8444
rect -936 -8508 -935 -8444
rect -1137 -8509 -935 -8508
rect -1137 -9991 -1061 -8509
rect 344 -9217 420 -7735
rect 2963 -8469 3410 -8468
rect 2963 -8533 3269 -8469
rect 3409 -8533 3410 -8469
rect 2963 -8534 3410 -8533
rect 2963 -8723 3039 -8534
rect 2495 -8789 3039 -8723
rect 344 -9218 546 -9217
rect 344 -9282 345 -9218
rect 545 -9282 546 -9218
rect 344 -9283 546 -9282
rect -1137 -9992 -935 -9991
rect -1137 -10056 -1136 -9992
rect -936 -10056 -935 -9992
rect -1137 -10057 -935 -10056
rect -1137 -10264 -1061 -10057
rect 344 -10264 420 -9283
rect 2495 -9369 2571 -8789
rect 2963 -8984 3039 -8789
rect 2963 -8985 3410 -8984
rect 2963 -9049 3269 -8985
rect 3409 -9049 3410 -8985
rect 2963 -9050 3410 -9049
rect 1965 -9370 2571 -9369
rect 1965 -9444 1966 -9370
rect 2566 -9444 2571 -9370
rect 1965 -9445 2571 -9444
rect 3144 -9277 3217 -9239
rect -1137 -10340 420 -10264
rect 3144 -9636 3149 -9277
rect 3214 -9636 3217 -9277
rect 3144 -9731 3217 -9636
rect 3144 -10090 3149 -9731
rect 3214 -10090 3217 -9731
rect -406 -10452 -329 -10340
rect 3144 -10452 3217 -10090
rect -406 -10528 3217 -10452
<< labels >>
rlabel metal2 14185 -1227 14185 -1227 3 vo3
port 1 e
rlabel metal3 -6150 -956 -6150 -956 5 vin_p
port 2 s
rlabel metal3 -8592 -989 -8592 -989 5 vin_n
port 3 s
rlabel metal4 895 7673 895 7673 3 vcc
port 4 e
rlabel metal4 -10692 -78 -10692 -78 7 vss
port 5 w
rlabel metal2 -1902 7526 -1902 7526 7 2nd_3_OTA_0.vcc
rlabel metal2 -1806 -1900 -1806 -1900 7 2nd_3_OTA_0.vss
rlabel metal1 -2007 3812 -2007 3812 7 2nd_3_OTA_0.vd1
rlabel metal1 -2008 3497 -2008 3497 7 2nd_3_OTA_0.vd2
rlabel metal4 7148 -1092 7148 -1092 7 2nd_3_OTA_0.vd4
rlabel metal3 7147 -1280 7147 -1280 7 2nd_3_OTA_0.vd3
rlabel metal2 6793 -1955 6793 -1955 5 2nd_3_OTA_0.vb1
rlabel metal2 3891 -10406 3891 -10406 5 OTA_vref_0.vcc
rlabel metal2 -1468 -10374 -1468 -10374 5 OTA_vref_0.vss
rlabel metal2 3005 -2773 3005 -2773 1 OTA_vref_0.vb
rlabel metal4 4081 -6638 4081 -6638 3 OTA_vref_0.vb1
rlabel metal2 3787 -7943 3787 -7943 1 OTA_vref_0.OTA_vref_stage2_0.vcc
rlabel metal2 2196 -8417 2196 -8417 1 OTA_vref_0.OTA_vref_stage2_0.vss
rlabel metal2 2516 -8448 2516 -8448 1 OTA_vref_0.OTA_vref_stage2_0.vref0
rlabel metal1 3196 -8015 3196 -8015 1 OTA_vref_0.OTA_vref_stage2_0.vr
rlabel metal2 3005 -2777 3005 -2777 1 OTA_vref_0.OTA_vref_stage2_0.vb
rlabel metal4 4073 -6642 4073 -6642 3 OTA_vref_0.OTA_vref_stage2_0.vb1
rlabel metal2 3890 -10392 3890 -10392 5 OTA_vref_0.OTA_vref_stage1_0.vcc
rlabel metal2 -1474 -10364 -1474 -10364 5 OTA_vref_0.OTA_vref_stage1_0.vss
rlabel metal3 1830 -8921 1830 -8921 3 OTA_vref_0.OTA_vref_stage1_0.vref0
rlabel metal1 3192 -8328 3192 -8328 1 OTA_vref_0.OTA_vref_stage1_0.vr
flabel locali 2206 -9753 2310 -9505 0 FreeSans 400 0 0 0 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter
flabel locali 1635 -9694 1684 -9593 0 FreeSans 400 0 0 0 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Collector
flabel locali 1794 -9717 1834 -9599 0 FreeSans 400 0 0 0 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Base
rlabel metal3 -6145 -400 -6145 -400 5 OTA_stage1_0.vin_p
rlabel metal3 -8611 -404 -8611 -404 5 OTA_stage1_0.vin_n
rlabel metal3 -9378 -406 -9378 -406 5 OTA_stage1_0.vb
rlabel metal2 -10396 5628 -10396 5628 7 OTA_stage1_0.vcc
rlabel metal2 -10398 -108 -10398 -108 7 OTA_stage1_0.vss
rlabel metal1 -2223 3813 -2223 3813 3 OTA_stage1_0.vd1
rlabel metal1 -2222 3501 -2222 3501 3 OTA_stage1_0.vd2
rlabel metal2 12164 2611 12164 2611 3 3rd_3_OTA_0.vcc
rlabel metal2 8412 -3643 8412 -3643 7 3rd_3_OTA_0.vss
rlabel metal2 12727 -1213 12727 -1213 3 3rd_3_OTA_0.vo3
rlabel metal1 7883 -1275 7883 -1275 7 3rd_3_OTA_0.vd3
rlabel metal1 7883 -1098 7883 -1098 7 3rd_3_OTA_0.vd4
rlabel metal3 10568 -3974 10568 -3974 7 3rd_3_OTA_0.vd1
rlabel metal3 8170 -2736 8170 -2736 7 3rd_3_OTA_0.vb
<< end >>
