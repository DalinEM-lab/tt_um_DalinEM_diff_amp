magic
tech sky130A
magscale 1 2
timestamp 1737772033
<< metal1 >>
rect 25795 5219 26678 5229
rect 25795 5129 26508 5219
rect 26498 4893 26508 5129
rect 26668 4893 26678 5219
<< via1 >>
rect 26508 4893 26668 5219
<< metal2 >>
rect 25822 7165 26855 7175
rect 25822 6786 26073 7165
rect 25822 6776 26855 6786
rect 25822 6775 26222 6776
rect 26508 5219 26668 5229
rect 26508 4883 26668 4893
rect 13344 1493 17814 1503
rect 14082 1113 17814 1493
rect 13344 1103 17814 1113
<< via2 >>
rect 26073 6786 26855 7165
rect 26508 4893 26668 5219
rect 13344 1113 14082 1493
<< metal3 >>
rect 26063 6776 26073 7174
rect 26855 6776 26865 7174
rect 26498 5219 26678 5224
rect 26498 4893 26508 5219
rect 26668 4893 26678 5219
rect 26498 4888 26678 4893
rect 13334 1104 13344 1502
rect 14083 1104 14093 1502
rect 18743 1028 18923 1029
rect 14906 1027 18923 1028
rect 14906 849 14930 1027
rect 15412 849 18923 1027
rect 14906 848 18923 849
rect 19516 782 19696 1047
rect 19168 604 19178 782
rect 19660 604 19696 782
rect 19516 603 19696 604
rect 21974 782 22154 1002
rect 21974 604 22018 782
rect 22500 604 22510 782
rect 21974 603 22154 604
<< via3 >>
rect 26073 7165 26855 7174
rect 26073 6786 26855 7165
rect 26073 6776 26855 6786
rect 26508 4893 26668 5219
rect 13344 1493 14083 1502
rect 13344 1113 14082 1493
rect 14082 1113 14083 1493
rect 13344 1104 14083 1113
rect 14930 849 15412 1027
rect 19178 604 19660 782
rect 22018 604 22500 782
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 14414 44152 14474 45152
rect 14966 44152 15026 45152
rect 15518 44152 15578 45152
rect 16070 44152 16130 45152
rect 16622 44152 16682 45152
rect 17174 44152 17234 45152
rect 17726 44152 17786 45152
rect 18278 44152 18338 45152
rect 18830 44152 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 400 43752 18890 44152
rect 400 1503 800 43752
rect 31400 7175 31800 44152
rect 25981 7174 31800 7175
rect 25981 6776 26073 7174
rect 26855 6776 31800 7174
rect 25981 6775 31800 6776
rect 26498 5219 26678 5229
rect 26498 4893 26508 5219
rect 26668 4893 26678 5219
rect 400 1502 14084 1503
rect 400 1104 13344 1502
rect 14083 1104 14084 1502
rect 400 1103 14084 1104
rect 400 1000 800 1103
rect 14906 1027 15413 1028
rect 14906 849 14930 1027
rect 15412 849 15413 1027
rect 14906 848 15413 849
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 848
rect 18770 782 19696 783
rect 18770 604 19178 782
rect 19660 604 19696 782
rect 18770 603 19696 604
rect 21974 782 22814 783
rect 21974 604 22018 782
rect 22500 604 22814 782
rect 21974 603 22814 604
rect 18770 0 18950 603
rect 22634 0 22814 603
rect 26498 0 26678 4893
rect 31400 1000 31800 6775
rect 30362 0 30542 200
use diff_final_v0  diff_final_v0_0 ~/Dalin/Projects/tinytape/diff_files
timestamp 1737769985
transform 1 0 6811 0 1 3794
box 10993 -2832 19171 3381
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 31400 1000 31800 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 1000 800 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
