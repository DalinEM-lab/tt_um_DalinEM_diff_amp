magic
tech sky130A
magscale 1 2
timestamp 1740775395
<< metal1 >>
rect -237 5771 0 5871
rect -257 5586 98 5686
rect 0 5462 98 5586
<< metal2 >>
rect 422 9631 2594 9641
rect 422 9451 2594 9461
rect -469 7417 319 7818
rect 69 2617 366 2627
rect -8486 1744 -8253 2145
rect -2133 1526 -1367 1845
rect 69 1840 366 1850
rect -7472 1495 -7292 1505
rect -7292 1394 -2999 1494
rect -7472 1384 -7292 1394
rect -3099 -1395 -2999 1394
rect -2133 1439 381 1526
rect -1469 977 381 1439
rect -2133 967 -1469 977
rect 8766 -199 8845 59
rect 8679 -209 8845 -199
rect -939 -406 -371 -266
rect 8679 -319 8845 -309
rect -939 -416 -365 -406
rect -939 -725 -365 -715
rect -3099 -1495 -1097 -1395
rect -2133 -2122 -1470 -2112
rect -1470 -2335 -833 -2122
rect -2133 -2345 -1470 -2335
rect -2133 -5819 -1469 -5809
rect -1469 -6016 -80 -5820
rect -2133 -6026 -1469 -6016
<< via2 >>
rect 422 9461 2594 9631
rect 69 1850 366 2617
rect -7472 1394 -7292 1495
rect -2133 977 -1469 1439
rect 8679 -309 8845 -209
rect -939 -715 -365 -416
rect -2133 -2335 -1470 -2122
rect -2133 -6016 -1469 -5819
<< metal3 >>
rect 412 9631 2604 9636
rect 412 9461 422 9631
rect 2594 9461 2604 9631
rect 412 9456 2604 9461
rect 59 2617 376 2622
rect 59 1850 69 2617
rect 366 1850 376 2617
rect 59 1845 376 1850
rect -7472 1500 -7292 1660
rect -7482 1495 -7282 1500
rect -7482 1394 -7472 1495
rect -7292 1394 -7282 1495
rect -7482 1389 -7282 1394
rect -6699 1320 -6519 1640
rect -4241 1298 -4061 1657
rect -2143 1439 -1459 1444
rect -2143 977 -2133 1439
rect -1469 977 -1459 1439
rect -2143 972 -1459 977
rect 8669 -209 8855 -204
rect 8669 -309 8679 -209
rect 8845 -309 8855 -209
rect 8669 -314 8855 -309
rect -949 -416 -355 -411
rect -949 -715 -939 -416
rect -365 -715 -355 -416
rect -949 -720 -355 -715
rect -2143 -2122 -1460 -2117
rect -2143 -2335 -2133 -2122
rect -1470 -2335 -1460 -2122
rect -2143 -2340 -1460 -2335
rect -2143 -5819 -1459 -5814
rect -2143 -6016 -2133 -5819
rect -1469 -6016 -1459 -5819
rect -2143 -6021 -1459 -6016
<< via3 >>
rect 422 9461 2594 9631
rect 69 1850 366 2617
rect -2133 977 -1469 1439
rect 8679 -309 8845 -209
rect -939 -715 -365 -416
rect -2133 -2335 -1470 -2122
rect -2133 -6016 -1469 -5819
<< metal4 >>
rect 156 9631 2794 9928
rect 156 9461 422 9631
rect 2594 9461 2794 9631
rect 156 9423 2794 9461
rect 68 2617 367 2618
rect -940 1850 69 2617
rect 366 1850 367 2617
rect -940 1849 -377 1850
rect 68 1849 367 1850
rect -2134 1439 -1468 1440
rect -2134 977 -2133 1439
rect -1469 977 -1468 1439
rect -2134 976 -1468 977
rect -2133 -2121 -1469 976
rect -939 -415 -377 1849
rect 8987 820 9167 1000
rect 8678 -209 8846 -208
rect 2718 -309 8679 -209
rect 8845 -309 8846 -209
rect 2718 -370 2784 -309
rect 8678 -310 8846 -309
rect -940 -416 -364 -415
rect -940 -715 -939 -416
rect -365 -715 -364 -416
rect -940 -716 -364 -715
rect -2134 -2122 -1469 -2121
rect -2134 -2335 -2133 -2122
rect -1470 -2335 -1469 -2122
rect -2134 -2336 -1469 -2335
rect -2133 -5818 -1469 -2336
rect -2134 -5819 -1468 -5818
rect -2134 -6016 -2133 -5819
rect -1469 -6016 -1468 -5819
rect -2134 -6017 -1468 -6016
use OTA_stage1  OTA_stage1_0 ~/Project_tinytape/magic/mag/OTA_stage1
timestamp 1740520188
transform 1 0 -19404 0 1 4436
box 10993 -2832 19171 3381
use OTA_stage2  OTA_stage2_0 ~/Project_tinytape/magic/mag/OTA_stage2
timestamp 1740515472
transform 1 0 -6296 0 1 5137
box 6296 -5137 15627 4514
use OTA_vref  OTA_vref_0 ~/Project_tinytape/magic/mag/OTA_vref
timestamp 1740539468
transform -1 0 6640 0 -1 -436
box 0 -73 7756 5648
<< labels >>
rlabel metal2 -8477 1929 -8477 1929 7 vss
port 1 w
rlabel metal4 2791 9774 2791 9774 3 vcc
port 2 e
rlabel metal4 9166 905 9166 905 3 vo
port 3 e
rlabel metal3 -4161 1299 -4161 1299 5 vin_p
port 4 s
rlabel metal3 -6618 1321 -6618 1321 5 vin_n
port 5 s
<< end >>
