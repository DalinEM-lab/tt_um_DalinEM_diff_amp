* NGSPICE file created from 2_OTA_flat.ext - technology: sky130A

.subckt x2_OTA_flat vss vcc vo vin_p vin_n
X0 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 a_n27_n4200.t47 vss.t65 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X1 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 OTA_vref_0.OTA_vref_stage2_0.vr.t19 vss.t42 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X2 OTA_vref_0.OTA_vref_stage2_0.vr.t18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 vss.t40 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X3 a_n832_n2063# a_n832_n2063# OTA_vref_0.vb vss.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=11600,516 d=5800,258
X4 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 a_n27_n4200.t45 vss.t64 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X5 a_n8089_3635# vin_p.t0 OTA_stage2_0.vd2.t0 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X6 OTA_vref_0.OTA_vref_stage2_0.vr.t17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 vss.t36 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X7 a_2980_n1975# a_3038_n2063# a_3038_n2063# vss.t78 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X8 a_458_n2063# a_458_n2063# a_400_n1975# vss.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X9 a_2980_n1975# a_1748_n2063# OTA_vref_0.vb1.t4 vss.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X10 a_400_n1975# a_458_n2063# a_458_n2063# vss.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X11 a_959_2177.t3 OTA_stage2_0.vd1.t5 vo.t1 vcc.t21 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X12 OTA_vref_0.vb1.t3 a_1748_n2063# a_1748_n2063# vss.t8 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X13 OTA_vref_0.vb1.t5 a_458_n2063# a_400_n1975# vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X14 a_959_2177.t2 OTA_stage2_0.vd1.t6 vo.t3 vcc.t20 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X15 vcc.t17 OTA_vref_0.OTA_vref_stage2_0.vr.t20 a_458_n2063# vcc.t16 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X16 vcc.t15 OTA_vref_0.OTA_vref_stage2_0.vr.t21 OTA_vref_0.vb vcc.t14 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X17 a_400_n1975# a_458_n2063# a_458_n2063# vss.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X18 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 a_n27_n4200.t46 vss.t63 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X19 OTA_vref_0.OTA_vref_stage2_0.vr.t16 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X20 vss.t67 a_521_2177.t12 vo.t6 vss.t66 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X21 vss.t72 a_521_2177.t13 vo.t7 vss.t71 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X22 a_521_2177.t11 OTA_stage2_0.vd2.t3 a_959_2177.t6 vcc.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X23 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 OTA_vref_0.OTA_vref_stage2_0.vr.t15 vss.t34 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X24 OTA_vref_0.OTA_vref_stage2_0.vr.t14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 vss.t46 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X25 vcc.t27 OTA_stage2_0.vd2.t0 OTA_stage2_0.vd2.t1 vcc.t25 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X26 a_521_2177.t7 a_521_2177.t6 vss.t3 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X27 OTA_vref_0.OTA_vref_stage2_0.vref0.t0 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 OTA_vref_0.OTA_vref_stage2_0.vr.t13 vss.t44 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X28 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 OTA_vref_0.OTA_vref_stage2_0.vr.t12 vss.t30 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X29 a_959_2177.t10 OTA_vref_0.vb1.t6 vcc.t35 vcc.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X30 a_n27_n4200.t44 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 vss.t59 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X31 a_8294_3178.t1 OTA_stage2_0.vd1.t2 sky130_fd_pr__cap_mim_m3_1 l=20 w=20
X32 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 OTA_vref_0.OTA_vref_stage2_0.vr.t11 vss.t38 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X33 vcc.t33 OTA_vref_0.vb1.t7 a_959_2177.t8 vcc.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=81200,2916 d=40600,1458
X34 vss.t57 a_n27_n4200.t26 a_n27_n4200.t27 vss.t56 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X35 vo.t8 a_521_2177.t14 vss.t79 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X36 a_n27_n4200.t38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 vss.t62 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X37 a_n27_n4200.t39 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 vss.t65 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X38 a_n27_n4200.t40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 vss.t64 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X39 vcc.t26 OTA_stage2_0.vd2.t0 OTA_stage2_0.vd1.t3 vcc.t25 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=20880,836 d=10440,418
X40 a_n27_n4200.t41 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 vss.t61 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X41 a_521_2177.t10 OTA_stage2_0.vd2.t4 a_959_2177.t4 vcc.t18 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X42 a_2980_n1975# a_3038_n2063# a_3038_n2063# vss.t77 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X43 OTA_vref_0.OTA_vref_stage2_0.vr.t10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 vss.t32 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X44 a_959_2177.t11 OTA_vref_0.vb1.t8 vcc.t31 vcc.t30 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=81200,2916
X45 a_n27_n4200.t42 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 vss.t60 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X46 OTA_stage2_0.vd1.t4 OTA_stage2_0.vd2.t0 vcc.t24 vcc.t22 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X47 a_3038_n2063# a_3038_n2063# a_2980_n1975# vss.t76 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X48 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 OTA_vref_0.OTA_vref_stage2_0.vr.t9 vss.t28 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X49 vcc.t29 OTA_vref_0.vb1.t9 a_959_2177.t9 vcc.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=7 l=1.8
**devattr s=40600,1458 d=40600,1458
X50 vss.t55 a_n27_n4200.t2 a_n27_n4200.t3 vss.t54 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X51 a_959_2177.t5 OTA_stage2_0.vd2.t5 a_521_2177.t9 vcc.t21 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X52 a_n27_n4200.t43 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 vss.t63 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X53 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 OTA_vref_0.OTA_vref_stage2_0.vr.t8 vss.t26 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X54 vss.t53 a_n27_n4200.t28 a_n27_n4200.t29 vss.t52 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X55 a_n27_n4200.t32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 vss.t58 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X56 vss.t51 a_n27_n4200.t4 a_n27_n4200.t5 vss.t50 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X57 a_n27_n4200.t7 a_n27_n4200.t6 vss.t49 vss.t48 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X58 a_400_n1975# a_n832_n2063# OTA_vref_0.vb vss.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=5800,258 d=5800,258
X59 vcc.t13 OTA_vref_0.OTA_vref_stage2_0.vr.t22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 vcc.t12 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=11600,516 d=5800,258
X60 vss.t47 a_n27_n4200.t30 a_n27_n4200.t31 vss.t46 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X61 a_n27_n4200.t19 a_n27_n4200.t18 vss.t45 vss.t44 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X62 OTA_stage2_0.vd2.t0 vin_p.t1 a_n8089_3635# vss.t12 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X63 a_n27_n4200.t15 a_n27_n4200.t14 vss.t43 vss.t42 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X64 vss.t41 a_n27_n4200.t20 a_n27_n4200.t21 vss.t40 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X65 a_n27_n4200.t9 a_n27_n4200.t8 vss.t39 vss.t38 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X66 vss.t70 a_521_2177.t4 a_521_2177.t5 vss.t66 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X67 vss.t37 a_n27_n4200.t22 a_n27_n4200.t23 vss.t36 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X68 a_1748_n2063# a_1748_n2063# OTA_vref_0.vb1.t2 vss.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X69 a_959_2177.t7 OTA_stage2_0.vd2.t6 a_521_2177.t8 vcc.t20 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=174000,6116 d=87000,3058
X70 OTA_stage2_0.vd2.t2 OTA_stage2_0.vd2.t0 vcc.t23 vcc.t22 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.8 l=18
**devattr s=10440,418 d=20880,836
X71 OTA_vref_0.vb a_n832_n2063# a_n832_n2063# vss.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X72 OTA_stage2_0.vd1.t1 vin_n.t0 a_n8089_3635# vss.t69 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.966667 ps=7.053333 w=6 l=12
**devattr s=34800,1258 d=69600,2516
X73 OTA_vref_0.vb a_n832_n2063# a_n832_n2063# vss.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.548 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X74 vss.t73 a_521_2177.t2 a_521_2177.t3 vss.t71 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=17400,716 d=8700,358
X75 vss.t63 vss.t68 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X76 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 a_n27_n4200.t37 vss.t62 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X77 a_n832_n2063# a_n832_n2063# OTA_vref_0.vb vss.t21 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.174 ps=1.548 w=1 l=1
**devattr s=5800,258 d=5800,258
X78 a_3038_n2063# a_3038_n2063# a_2980_n1975# vss.t75 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X79 vo.t4 OTA_stage2_0.vd1.t7 a_959_2177.t1 vcc.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=87000,3058
X80 vo.t0 a_521_2177.t15 vss.t2 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=8700,358
X81 a_8294_3178.t0 vo.t5 vss.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1
X82 a_458_n2063# a_458_n2063# a_400_n1975# vss.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X83 a_1748_n2063# a_1748_n2063# OTA_vref_0.vb1.t1 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=5800,258
X84 a_n27_n4200.t13 a_n27_n4200.t12 vss.t35 vss.t34 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X85 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 a_n27_n4200.t33 vss.t61 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X86 vcc.t11 OTA_vref_0.OTA_vref_stage2_0.vr.t23 a_n832_n2063# vcc.t10 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X87 vss.t33 a_n27_n4200.t24 a_n27_n4200.t25 vss.t32 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=46400,1716
X88 OTA_vref_0.vb1.t0 a_1748_n2063# a_1748_n2063# vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X89 vcc.t7 OTA_vref_0.OTA_vref_stage2_0.vr.t0 OTA_vref_0.OTA_vref_stage2_0.vr.t1 vcc.t6 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=5800,316 d=2900,158
X90 vcc.t9 OTA_vref_0.OTA_vref_stage2_0.vr.t24 a_3038_n2063# vcc.t8 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X91 a_n27_n4200.t17 a_n27_n4200.t16 vss.t31 vss.t30 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X92 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 a_n27_n4200.t34 vss.t60 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X93 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 a_n27_n4200.t35 vss.t59 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 OTA_vref_0.OTA_vref_stage2_0.vr.t25 vcc.t5 vcc.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=1
**devattr s=5800,258 d=11600,516
X95 a_521_2177.t1 a_521_2177.t0 vss.t11 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1.5 l=9.4
**devattr s=8700,358 d=17400,716
X96 vo.t2 OTA_stage2_0.vd1.t8 a_959_2177.t0 vcc.t18 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=15 l=1.9
**devattr s=87000,3058 d=174000,6116
X97 a_n27_n4200.t1 a_n27_n4200.t0 vss.t29 vss.t28 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X98 OTA_vref_0.OTA_vref_stage2_0.vref0.t32 a_3038_n2063# a_2980_n1975# vss.t74 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=11600,516
X99 vcc.t3 OTA_vref_0.OTA_vref_stage2_0.vr.t26 a_1748_n2063# vcc.t2 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=11600,516
X100 OTA_vref_0.OTA_vref_stage2_0.vr.t7 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 vss.t54 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X101 a_n8089_3635# vin_n.t1 OTA_stage2_0.vd1.t0 vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.966667 pd=7.053333 as=0 ps=0 w=6 l=12
**devattr s=69600,2516 d=34800,1258
X102 OTA_vref_0.OTA_vref_stage2_0.vr.t6 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 vss.t56 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X103 a_n8089_3635# OTA_vref_0.vb vss.t14 vss.t13 sky130_fd_pr__nfet_01v8 ad=0.483333 pd=3.526667 as=0 ps=0 w=3 l=5
**devattr s=34800,1316 d=34800,1316
X104 a_n27_n4200.t11 a_n27_n4200.t10 vss.t27 vss.t26 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=23200,858
X105 OTA_vref_0.OTA_vref_stage2_0.vr.t5 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 vss.t50 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X106 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 a_n27_n4200.t36 vss.t58 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X107 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 OTA_vref_0.OTA_vref_stage2_0.vr.t4 vss.t48 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=23200,858 d=23200,858
X108 OTA_vref_0.OTA_vref_stage2_0.vr.t3 OTA_vref_0.OTA_vref_stage2_0.vr.t2 vcc.t1 vcc.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=0.5 l=2
**devattr s=2900,158 d=5800,316
R0 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 1594.54
R1 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 235.982
R2 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 235.978
R3 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 190.305
R4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 190.305
R5 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 190.305
R6 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 190.305
R7 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 190.305
R8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 190.305
R9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 190.305
R10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 190.305
R11 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 190.305
R12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 190.305
R13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 190.305
R14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 190.305
R15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 95.392
R16 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 95.3648
R17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 95.1871
R18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 95.1789
R19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 95.1789
R20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 95.1754
R21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 95.1707
R22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 95.1542
R23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 95.1542
R24 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 94.8314
R25 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 94.8314
R26 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 94.8314
R27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 94.8314
R28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 94.8314
R29 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 94.8314
R30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 94.8314
R31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 94.8314
R32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 94.8314
R33 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 94.8314
R34 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 94.8314
R35 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 94.8314
R36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 94.8314
R37 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 94.8314
R38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 94.8314
R39 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 94.8314
R40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 94.8314
R41 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 84.0884
R42 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 83.5719
R43 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 83.5719
R44 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 83.5719
R45 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 83.5719
R46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 73.19
R47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 26.074
R48 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 26.074
R49 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 26.074
R50 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 25.7843
R51 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 10.2822
R52 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 9.66384
R53 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 7.22993
R54 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 7.22993
R55 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 7.22819
R56 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 6.83022
R57 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 6.81633
R58 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 6.81633
R59 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 6.81633
R60 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 6.75312
R61 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 2.36206
R62 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 2.29815
R63 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 1.86108
R64 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 1.86108
R65 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 1.86108
R66 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 1.86108
R67 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 1.86108
R68 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 1.86108
R69 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 1.86108
R70 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 1.55316
R71 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 1.5505
R72 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 1.5505
R73 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 1.5505
R74 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 1.5505
R75 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 1.28702
R76 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 1.25468
R77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 1.14402
R78 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 1.1424
R79 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 1.11251
R80 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 1.10979
R81 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 1.10164
R82 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 1.10164
R83 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 1.09892
R84 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 1.08805
R85 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 1.08262
R86 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 1.07024
R87 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 1.06903
R88 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 1.06903
R89 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 1.0237
R90 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.885803
R91 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 0.77514
R92 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 0.756696
R93 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 0.701365
R94 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 0.645119
R95 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 0.645119
R96 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n66 0.645119
R97 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 0.645119
R98 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n57 0.645119
R99 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 0.645119
R100 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 0.645119
R101 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n47 0.645119
R102 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 0.645119
R103 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 0.645119
R104 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 0.645119
R105 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n38 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 0.645119
R106 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 0.645119
R107 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 0.645119
R108 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 0.645119
R109 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n28 0.645119
R110 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 0.645119
R111 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 0.645119
R112 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n17 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 0.645119
R113 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n19 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 0.645119
R114 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 0.645119
R115 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 0.645119
R116 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n9 0.645119
R117 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 0.645117
R118 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 0.590702
R119 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 0.495065
R120 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 0.495065
R121 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 0.481478
R122 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 0.481478
R123 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 0.475521
R124 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 0.470609
R125 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 0.470609
R126 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 0.465174
R127 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 0.465174
R128 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 0.465174
R129 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 0.459844
R130 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 0.459739
R131 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 0.459739
R132 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 0.446152
R133 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 0.446152
R134 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 0.445943
R135 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 0.443435
R136 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 0.440717
R137 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 0.440717
R138 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 0.434551
R139 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 0.431769
R140 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 0.414484
R141 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 0.410839
R142 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 0.410839
R143 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.408265
R144 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 0.408265
R145 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.408265
R146 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 0.408265
R147 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.407145
R148 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 0.407145
R149 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 0.405635
R150 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 0.405635
R151 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 0.290206
R152 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 0.203382
R153 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 0.0209918
R154 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 0.0209918
R155 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 0.0209918
R156 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 0.0209918
R157 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 0.0183279
R158 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 0.0074695
R159 a_n27_n4200.n1 a_n27_n4200.t22 94.9536
R160 a_n27_n4200.n1 a_n27_n4200.n0 0.400892
R161 a_n27_n4200.n33 a_n27_n4200.t16 190.305
R162 a_n27_n4200.t16 a_n27_n4200.n9 190.305
R163 a_n27_n4200.n33 a_n27_n4200.n8 0.559233
R164 a_n27_n4200.t4 a_n27_n4200.n8 94.8744
R165 a_n27_n4200.n30 a_n27_n4200.n19 0.302364
R166 a_n27_n4200.n19 a_n27_n4200.t26 95.0028
R167 a_n27_n4200.t18 a_n27_n4200.n29 94.9085
R168 a_n27_n4200.n34 a_n27_n4200.t6 190.305
R169 a_n27_n4200.t6 a_n27_n4200.n12 190.305
R170 a_n27_n4200.n34 a_n27_n4200.n13 0.561351
R171 a_n27_n4200.t20 a_n27_n4200.n13 94.8733
R172 a_n27_n4200.n5 a_n27_n4200.t28 94.8439
R173 a_n27_n4200.n5 a_n27_n4200.n4 0.620271
R174 a_n27_n4200.n6 a_n27_n4200.t8 190.305
R175 a_n27_n4200.t8 a_n27_n4200.n4 190.305
R176 a_n27_n4200.t2 a_n27_n4200.n3 94.9565
R177 a_n27_n4200.n2 a_n27_n4200.n3 0.39509
R178 a_n27_n4200.n16 a_n27_n4200.t30 190.305
R179 a_n27_n4200.n14 a_n27_n4200.t30 190.305
R180 a_n27_n4200.n15 a_n27_n4200.t0 94.8665
R181 a_n27_n4200.n15 a_n27_n4200.n14 0.574949
R182 a_n27_n4200.n48 a_n27_n4200.t10 95.1811
R183 a_n27_n4200.n37 a_n27_n4200.t24 95.1783
R184 a_n27_n4200.n22 a_n27_n4200.n38 22.3176
R185 a_n27_n4200.n24 a_n27_n4200.n43 22.2301
R186 a_n27_n4200.n25 a_n27_n4200.n49 22.2284
R187 a_n27_n4200.n26 a_n27_n4200.n50 22.2284
R188 a_n27_n4200.n26 a_n27_n4200.n44 22.2284
R189 a_n27_n4200.n24 a_n27_n4200.n42 22.2284
R190 a_n27_n4200.n27 a_n27_n4200.n41 22.2284
R191 a_n27_n4200.n28 a_n27_n4200.n36 22.2284
R192 a_n27_n4200.n57 a_n27_n4200.n27 22.2284
R193 a_n27_n4200.n21 a_n27_n4200.n47 22.1884
R194 a_n27_n4200.n21 a_n27_n4200.n46 22.1884
R195 a_n27_n4200.n20 a_n27_n4200.n45 22.1884
R196 a_n27_n4200.n20 a_n27_n4200.n53 22.1884
R197 a_n27_n4200.n23 a_n27_n4200.n54 22.1884
R198 a_n27_n4200.n23 a_n27_n4200.n40 22.1884
R199 a_n27_n4200.n22 a_n27_n4200.n39 22.1884
R200 a_n27_n4200.n31 a_n27_n4200.n37 11.5566
R201 a_n27_n4200.n48 a_n27_n4200.n32 10.9335
R202 a_n27_n4200.n9 a_n27_n4200.n32 9.80925
R203 a_n27_n4200.n12 a_n27_n4200.n52 9.80925
R204 a_n27_n4200.n55 a_n27_n4200.n2 9.80925
R205 a_n27_n4200.n0 a_n27_n4200.n31 9.80925
R206 a_n27_n4200.n6 a_n27_n4200.n35 9.403
R207 a_n27_n4200.n51 a_n27_n4200.n30 9.39819
R208 a_n27_n4200.n16 a_n27_n4200.n56 9.39819
R209 a_n27_n4200.n37 a_n27_n4200.n28 4.9275
R210 a_n27_n4200.n25 a_n27_n4200.n48 4.79654
R211 a_n27_n4200.n22 a_n27_n4200.n0 2.24062
R212 a_n27_n4200.n23 a_n27_n4200.n2 2.23747
R213 a_n27_n4200.n20 a_n27_n4200.n11 1.89164
R214 a_n27_n4200.n12 a_n27_n4200.n11 0.719718
R215 a_n27_n4200.n10 a_n27_n4200.n21 1.88964
R216 a_n27_n4200.n10 a_n27_n4200.n9 0.723726
R217 a_n27_n4200.n17 a_n27_n4200.n16 0.692577
R218 a_n27_n4200.n17 a_n27_n4200.n27 1.90521
R219 a_n27_n4200.n7 a_n27_n4200.n24 1.87937
R220 a_n27_n4200.n7 a_n27_n4200.n6 0.744259
R221 a_n27_n4200.n26 a_n27_n4200.n18 1.94941
R222 a_n27_n4200.n49 a_n27_n4200.t37 4.3505
R223 a_n27_n4200.n49 a_n27_n4200.t11 4.3505
R224 a_n27_n4200.n50 a_n27_n4200.t27 4.3505
R225 a_n27_n4200.n50 a_n27_n4200.t39 4.3505
R226 a_n27_n4200.n44 a_n27_n4200.t33 4.3505
R227 a_n27_n4200.n44 a_n27_n4200.t19 4.3505
R228 a_n27_n4200.n43 a_n27_n4200.t29 4.3505
R229 a_n27_n4200.n43 a_n27_n4200.t44 4.3505
R230 a_n27_n4200.n42 a_n27_n4200.t36 4.3505
R231 a_n27_n4200.n42 a_n27_n4200.t9 4.3505
R232 a_n27_n4200.n41 a_n27_n4200.t31 4.3505
R233 a_n27_n4200.n41 a_n27_n4200.t40 4.3505
R234 a_n27_n4200.n36 a_n27_n4200.t25 4.3505
R235 a_n27_n4200.n36 a_n27_n4200.t43 4.3505
R236 a_n27_n4200.n47 a_n27_n4200.t5 4.3505
R237 a_n27_n4200.n47 a_n27_n4200.t38 4.3505
R238 a_n27_n4200.n46 a_n27_n4200.t47 4.3505
R239 a_n27_n4200.n46 a_n27_n4200.t17 4.3505
R240 a_n27_n4200.n45 a_n27_n4200.t21 4.3505
R241 a_n27_n4200.n45 a_n27_n4200.t41 4.3505
R242 a_n27_n4200.n53 a_n27_n4200.t35 4.3505
R243 a_n27_n4200.n53 a_n27_n4200.t7 4.3505
R244 a_n27_n4200.n54 a_n27_n4200.t3 4.3505
R245 a_n27_n4200.n54 a_n27_n4200.t32 4.3505
R246 a_n27_n4200.n40 a_n27_n4200.t45 4.3505
R247 a_n27_n4200.n40 a_n27_n4200.t13 4.3505
R248 a_n27_n4200.n39 a_n27_n4200.t23 4.3505
R249 a_n27_n4200.n39 a_n27_n4200.t42 4.3505
R250 a_n27_n4200.n38 a_n27_n4200.t46 4.3505
R251 a_n27_n4200.n38 a_n27_n4200.t15 4.3505
R252 a_n27_n4200.n57 a_n27_n4200.t34 4.3505
R253 a_n27_n4200.t1 a_n27_n4200.n57 4.3505
R254 a_n27_n4200.n25 a_n27_n4200.n21 2.55258
R255 a_n27_n4200.n23 a_n27_n4200.n22 2.02133
R256 a_n27_n4200.n56 a_n27_n4200.n31 1.86108
R257 a_n27_n4200.n56 a_n27_n4200.n55 1.86108
R258 a_n27_n4200.n55 a_n27_n4200.n35 1.86108
R259 a_n27_n4200.n52 a_n27_n4200.n35 1.86108
R260 a_n27_n4200.n52 a_n27_n4200.n51 1.86108
R261 a_n27_n4200.n51 a_n27_n4200.n32 1.86108
R262 a_n27_n4200.n26 a_n27_n4200.n25 1.74425
R263 a_n27_n4200.n10 a_n27_n4200.n33 1.38566
R264 a_n27_n4200.n34 a_n27_n4200.n11 1.38875
R265 a_n27_n4200.n18 a_n27_n4200.n29 1.67497
R266 a_n27_n4200.n27 a_n27_n4200.n28 1.613
R267 a_n27_n4200.n26 a_n27_n4200.n24 1.613
R268 a_n27_n4200.n23 a_n27_n4200.n20 1.613
R269 a_n27_n4200.n21 a_n27_n4200.n20 1.613
R270 a_n27_n4200.n19 a_n27_n4200.n18 0.302364
R271 a_n27_n4200.n6 a_n27_n4200.n5 0.620271
R272 a_n27_n4200.n16 a_n27_n4200.n15 0.574949
R273 a_n27_n4200.n13 a_n27_n4200.n12 0.561351
R274 a_n27_n4200.n9 a_n27_n4200.n8 0.559233
R275 a_n27_n4200.n24 a_n27_n4200.n27 1.0755
R276 a_n27_n4200.n30 a_n27_n4200.n29 0.491095
R277 a_n27_n4200.n4 a_n27_n4200.n7 1.50352
R278 a_n27_n4200.n17 a_n27_n4200.n14 1.39428
R279 a_n27_n4200.t12 a_n27_n4200.n3 95.226
R280 a_n27_n4200.t14 a_n27_n4200.n1 95.2318
R281 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.t32 88.7532
R282 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 22.2005
R283 OTA_vref_0.OTA_vref_stage2_0.vref0.n25 OTA_vref_0.OTA_vref_stage2_0.vref0.n24 21.8815
R284 OTA_vref_0.OTA_vref_stage2_0.vref0.n25 OTA_vref_0.OTA_vref_stage2_0.vref0.n23 21.5624
R285 OTA_vref_0.OTA_vref_stage2_0.vref0.n26 OTA_vref_0.OTA_vref_stage2_0.vref0.n22 21.5624
R286 OTA_vref_0.OTA_vref_stage2_0.vref0.n27 OTA_vref_0.OTA_vref_stage2_0.vref0.n21 21.5624
R287 OTA_vref_0.OTA_vref_stage2_0.vref0.n28 OTA_vref_0.OTA_vref_stage2_0.vref0.n20 21.5624
R288 OTA_vref_0.OTA_vref_stage2_0.vref0.n29 OTA_vref_0.OTA_vref_stage2_0.vref0.n19 21.5624
R289 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 21.5624
R290 OTA_vref_0.OTA_vref_stage2_0.vref0.n18 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 21.5603
R291 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 21.5445
R292 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 21.5445
R293 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 21.5445
R294 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 21.5445
R295 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 21.5445
R296 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 21.5445
R297 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 21.5445
R298 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 4.3505
R299 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 4.3505
R300 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 4.3505
R301 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 OTA_vref_0.OTA_vref_stage2_0.vref0.t0 4.3505
R302 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 4.3505
R303 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 4.3505
R304 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 4.3505
R305 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 4.3505
R306 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 4.3505
R307 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 4.3505
R308 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 4.3505
R309 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 4.3505
R310 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 4.3505
R311 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 4.3505
R312 OTA_vref_0.OTA_vref_stage2_0.vref0.n24 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 4.3505
R313 OTA_vref_0.OTA_vref_stage2_0.vref0.n24 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 4.3505
R314 OTA_vref_0.OTA_vref_stage2_0.vref0.n23 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 4.3505
R315 OTA_vref_0.OTA_vref_stage2_0.vref0.n23 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 4.3505
R316 OTA_vref_0.OTA_vref_stage2_0.vref0.n22 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 4.3505
R317 OTA_vref_0.OTA_vref_stage2_0.vref0.n22 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 4.3505
R318 OTA_vref_0.OTA_vref_stage2_0.vref0.n21 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 4.3505
R319 OTA_vref_0.OTA_vref_stage2_0.vref0.n21 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 4.3505
R320 OTA_vref_0.OTA_vref_stage2_0.vref0.n20 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 4.3505
R321 OTA_vref_0.OTA_vref_stage2_0.vref0.n20 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 4.3505
R322 OTA_vref_0.OTA_vref_stage2_0.vref0.n19 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 4.3505
R323 OTA_vref_0.OTA_vref_stage2_0.vref0.n19 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 4.3505
R324 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 4.3505
R325 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 4.3505
R326 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 4.3505
R327 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 4.3505
R328 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 4.3505
R329 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 4.3505
R330 OTA_vref_0.OTA_vref_stage2_0.vref0.n18 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 1.5282
R331 OTA_vref_0.OTA_vref_stage2_0.vref0.n28 OTA_vref_0.OTA_vref_stage2_0.vref0.n27 0.638711
R332 OTA_vref_0.OTA_vref_stage2_0.vref0.n26 OTA_vref_0.OTA_vref_stage2_0.vref0.n25 0.638711
R333 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 0.624699
R334 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 0.624699
R335 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 0.624699
R336 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n29 0.59171
R337 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 0.414842
R338 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 OTA_vref_0.OTA_vref_stage2_0.vref0.n18 0.366605
R339 OTA_vref_0.OTA_vref_stage2_0.vref0.n29 OTA_vref_0.OTA_vref_stage2_0.vref0.n28 0.319605
R340 OTA_vref_0.OTA_vref_stage2_0.vref0.n27 OTA_vref_0.OTA_vref_stage2_0.vref0.n26 0.319605
R341 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 0.296969
R342 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 0.296969
R343 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 0.296969
R344 vss.n280 vss.n279 3.00584e+06
R345 vss.n311 vss.n280 2.2308e+06
R346 vss.n311 vss.n310 1.408e+06
R347 vss.n382 vss.n381 50190.3
R348 vss.n381 vss.n380 43514.2
R349 vss.n292 vss.n284 27614.8
R350 vss.n306 vss.n284 27609
R351 vss.n292 vss.n285 27609
R352 vss.n306 vss.n285 27603.2
R353 vss.n313 vss.n98 26954.2
R354 vss.n313 vss.n277 26954.2
R355 vss.n315 vss.n98 26948.4
R356 vss.n315 vss.n277 26948.4
R357 vss.n20 vss.n5 25442
R358 vss.n20 vss.n6 25442
R359 vss.n11 vss.n5 25436.2
R360 vss.n11 vss.n6 25436.2
R361 vss.n381 vss.n22 25416
R362 vss.n361 vss.n47 17753.2
R363 vss.n361 vss.n48 17753.2
R364 vss.n363 vss.n47 17753.2
R365 vss.n363 vss.n48 17753.2
R366 vss.n307 vss.n22 7306.95
R367 vss.n107 vss.n102 7296
R368 vss.n111 vss.n107 6735.47
R369 vss.n14 vss.n3 6275.03
R370 vss.n383 vss.n3 6275.03
R371 vss.n14 vss.n4 6275.03
R372 vss.n383 vss.n4 6275.03
R373 vss.n309 vss.n49 5636.95
R374 vss.n312 vss.n311 5636.95
R375 vss.n308 vss.n283 5430.16
R376 vss.n28 vss.n25 4403.53
R377 vss.n379 vss.n24 4403.53
R378 vss.n379 vss.n25 4403.53
R379 vss.n380 vss.n23 3337.68
R380 vss.n114 vss.t10 3239.87
R381 vss.n291 vss.t66 2286.68
R382 vss.n332 vss.n331 1945.46
R383 vss.t71 vss.n308 1669.14
R384 vss.n310 vss.n309 1614.22
R385 vss.n380 vss.t10 1536.63
R386 vss.t66 vss.n290 1492.06
R387 vss.n304 vss.n286 903.91
R388 vss.n358 vss.n357 884.182
R389 vss.n290 vss.n23 738.096
R390 vss.n280 vss.n23 609.524
R391 vss.n349 vss.n59 585
R392 vss.n113 vss.n59 585
R393 vss.n348 vss.n347 585
R394 vss.n151 vss.n62 585
R395 vss.n156 vss.n155 585
R396 vss.n161 vss.n160 585
R397 vss.n163 vss.n162 585
R398 vss.n176 vss.n175 585
R399 vss.n174 vss.n173 585
R400 vss.n170 vss.n169 585
R401 vss.n168 vss.n71 585
R402 vss.n342 vss.n69 585
R403 vss.n344 vss.n343 585
R404 vss.n345 vss.n344 585
R405 vss.n181 vss.n53 585
R406 vss.n185 vss.n184 585
R407 vss.n190 vss.n189 585
R408 vss.n192 vss.n191 585
R409 vss.n212 vss.n211 585
R410 vss.n210 vss.n209 585
R411 vss.n202 vss.n196 585
R412 vss.n204 vss.n203 585
R413 vss.n198 vss.n197 585
R414 vss.n353 vss.n54 585
R415 vss.n353 vss.n352 585
R416 vss.n353 vss.n52 585
R417 vss.n330 vss.n100 585
R418 vss.n331 vss.n330 585
R419 vss.n329 vss.n99 585
R420 vss.n257 vss.n101 585
R421 vss.n260 vss.n259 585
R422 vss.n261 vss.n260 585
R423 vss.n226 vss.n224 585
R424 vss.n262 vss.n226 585
R425 vss.n266 vss.n265 585
R426 vss.n265 vss.n264 585
R427 vss.n256 vss.n255 585
R428 vss.n263 vss.n256 585
R429 vss.n251 vss.n227 585
R430 vss.n233 vss.n227 585
R431 vss.n231 vss.n228 585
R432 vss.n234 vss.n231 585
R433 vss.n246 vss.n245 585
R434 vss.n245 vss.n244 585
R435 vss.n237 vss.n232 585
R436 vss.n243 vss.n232 585
R437 vss.n241 vss.n240 585
R438 vss.n242 vss.n241 585
R439 vss.n239 vss.n236 585
R440 vss.n236 vss.n235 585
R441 vss.n115 vss.n68 585
R442 vss.n117 vss.n116 585
R443 vss.n120 vss.n118 585
R444 vss.n118 vss.n110 585
R445 vss.n126 vss.n125 585
R446 vss.n127 vss.n126 585
R447 vss.n109 vss.n105 585
R448 vss.n128 vss.n109 585
R449 vss.n130 vss.n106 585
R450 vss.n130 vss.n129 585
R451 vss.n143 vss.n142 585
R452 vss.n142 vss.n141 585
R453 vss.n132 vss.n131 585
R454 vss.n140 vss.n131 585
R455 vss.n138 vss.n137 585
R456 vss.n139 vss.n138 585
R457 vss.n95 vss.n93 585
R458 vss.n97 vss.n95 585
R459 vss.n335 vss.n334 585
R460 vss.n334 vss.n333 585
R461 vss.n96 vss.n94 585
R462 vss.n332 vss.n96 585
R463 vss.n310 vss.t1 550.812
R464 vss.n21 vss.t69 535.15
R465 vss.n12 vss.t4 535.15
R466 vss.n309 vss.t71 482.603
R467 vss.n10 vss.t12 449.248
R468 vss.t0 vss.n10 448.884
R469 vss.n113 vss.t63 403.053
R470 vss.n28 vss.n27 338.354
R471 vss.n63 vss.t63 322.904
R472 vss.n114 vss.n113 319.084
R473 vss.n308 vss.n307 312.86
R474 vss.n19 vss.n7 307.036
R475 vss.n30 vss.n25 292.5
R476 vss.n25 vss.t20 292.5
R477 vss.n26 vss.n24 292.5
R478 vss.n276 vss.n45 287.481
R479 vss.n360 vss.n46 281.336
R480 vss.n360 vss.n359 281.243
R481 vss.t25 vss.n281 277.521
R482 vss.n356 vss.n355 264.301
R483 vss.n373 vss.n372 262.366
R484 vss.n352 vss.n59 259.416
R485 vss.n380 vss.n379 259.197
R486 vss.n340 vss.n72 258.334
R487 vss.n351 vss.n350 257.99
R488 vss.n8 vss.n7 256.805
R489 vss.n316 vss.n276 255.26
R490 vss.n346 vss.n345 254.34
R491 vss.n345 vss.n64 254.34
R492 vss.n345 vss.n65 254.34
R493 vss.n345 vss.n66 254.34
R494 vss.n345 vss.n67 254.34
R495 vss.n354 vss.n353 254.34
R496 vss.n353 vss.n58 254.34
R497 vss.n353 vss.n57 254.34
R498 vss.n353 vss.n56 254.34
R499 vss.n353 vss.n55 254.34
R500 vss.n328 vss.n327 254.34
R501 vss.n112 vss.n111 254.34
R502 vss.n27 vss.n24 253.208
R503 vss.n34 vss.n32 252.304
R504 vss.n344 vss.n68 249.663
R505 vss.t28 vss.t60 242.357
R506 vss.t21 vss.t23 241.893
R507 vss.t23 vss.t25 241.893
R508 vss.t1 vss.n280 236.508
R509 vss.n278 vss.t28 235.781
R510 vss.t22 vss.n282 226.892
R511 vss.n294 vss.n293 223.468
R512 vss.n384 vss.n2 216.017
R513 vss.n114 vss.n63 215.269
R514 vss.t78 vss.t54 213.556
R515 vss.t75 vss.t58 213.556
R516 vss.t77 vss.t38 213.556
R517 vss.t9 vss.t59 213.556
R518 vss.t8 vss.t48 213.556
R519 vss.t6 vss.t40 213.556
R520 vss.t5 vss.t61 213.556
R521 vss.t56 vss.t17 213.556
R522 vss.t65 vss.t16 213.556
R523 vss.t30 vss.t19 213.556
R524 vss.t24 vss.t26 212.828
R525 vss.t74 vss.t34 204.142
R526 vss.n326 vss.n325 200.388
R527 vss.n357 vss.n50 200.317
R528 vss.n236 vss.n52 197
R529 vss.n115 vss.n114 195.238
R530 vss.t50 vss.t18 195.044
R531 vss.n330 vss.n329 187.249
R532 vss.n238 vss.n81 185
R533 vss.t68 vss.n81 185
R534 vss.n230 vss.n229 185
R535 vss.n248 vss.n247 185
R536 vss.n250 vss.n249 185
R537 vss.n254 vss.n253 185
R538 vss.n252 vss.n225 185
R539 vss.n268 vss.n267 185
R540 vss.n258 vss.n86 185
R541 vss.t68 vss.n86 185
R542 vss.n103 vss.n91 185
R543 vss.n183 vss.n182 185
R544 vss.n188 vss.n187 185
R545 vss.n186 vss.n180 185
R546 vss.n195 vss.n194 185
R547 vss.n193 vss.n179 185
R548 vss.n208 vss.n207 185
R549 vss.n206 vss.n205 185
R550 vss.n201 vss.n200 185
R551 vss.n199 vss.n60 185
R552 vss.n152 vss.n61 185
R553 vss.n154 vss.n153 185
R554 vss.n159 vss.n158 185
R555 vss.n157 vss.n150 185
R556 vss.n166 vss.n165 185
R557 vss.n164 vss.n149 185
R558 vss.n172 vss.n171 185
R559 vss.n167 vss.n73 185
R560 vss.n341 vss.n340 185
R561 vss.n119 vss.n72 185
R562 vss.n122 vss.n121 185
R563 vss.n124 vss.n123 185
R564 vss.n147 vss.n146 185
R565 vss.n145 vss.n144 185
R566 vss.n133 vss.n108 185
R567 vss.n135 vss.n134 185
R568 vss.n136 vss.n92 185
R569 vss.n337 vss.n336 185
R570 vss.n9 vss.n8 184.031
R571 vss.n283 vss.t62 182.826
R572 vss.n19 vss.n18 177.084
R573 vss.n22 vss.n21 176.556
R574 vss.n197 vss.n54 175.546
R575 vss.n203 vss.n202 175.546
R576 vss.n211 vss.n210 175.546
R577 vss.n191 vss.n190 175.546
R578 vss.n184 vss.n53 175.546
R579 vss.n260 vss.n101 175.546
R580 vss.n260 vss.n226 175.546
R581 vss.n265 vss.n226 175.546
R582 vss.n265 vss.n256 175.546
R583 vss.n256 vss.n227 175.546
R584 vss.n231 vss.n227 175.546
R585 vss.n245 vss.n231 175.546
R586 vss.n245 vss.n232 175.546
R587 vss.n241 vss.n232 175.546
R588 vss.n241 vss.n236 175.546
R589 vss.n118 vss.n117 175.546
R590 vss.n126 vss.n118 175.546
R591 vss.n126 vss.n109 175.546
R592 vss.n130 vss.n109 175.546
R593 vss.n142 vss.n130 175.546
R594 vss.n142 vss.n131 175.546
R595 vss.n138 vss.n131 175.546
R596 vss.n138 vss.n95 175.546
R597 vss.n334 vss.n95 175.546
R598 vss.n334 vss.n96 175.546
R599 vss.n344 vss.n69 175.546
R600 vss.n169 vss.n168 175.546
R601 vss.n175 vss.n174 175.546
R602 vss.n162 vss.n161 175.546
R603 vss.n155 vss.n62 175.546
R604 vss.n347 vss.n59 175.546
R605 vss.n292 vss.n291 172.708
R606 vss.n295 vss.n287 169.446
R607 vss.n353 vss.t60 169.087
R608 vss.n13 vss.t13 167.053
R609 vss.n382 vss.t13 167.053
R610 vss.n182 vss.n81 163.333
R611 vss.n279 vss.t46 152.179
R612 vss.n314 vss.t52 150.524
R613 vss.n123 vss.n122 150
R614 vss.n146 vss.n145 150
R615 vss.n134 vss.n133 150
R616 vss.n337 vss.n92 150
R617 vss.n171 vss.n73 150
R618 vss.n165 vss.n164 150
R619 vss.n158 vss.n157 150
R620 vss.n153 vss.n152 150
R621 vss.n200 vss.n199 150
R622 vss.n207 vss.n206 150
R623 vss.n194 vss.n193 150
R624 vss.n187 vss.n186 150
R625 vss.n91 vss.n86 150
R626 vss.n267 vss.n86 150
R627 vss.n253 vss.n252 150
R628 vss.n249 vss.n248 150
R629 vss.n229 vss.n81 150
R630 vss.n324 vss.n104 137.462
R631 vss.n355 vss.n354 132.721
R632 vss.n13 vss.n12 132.691
R633 vss.n380 vss.t20 131.666
R634 vss.n116 vss.n115 129.202
R635 vss.n116 vss.n110 129.202
R636 vss.n127 vss.n110 129.202
R637 vss.n128 vss.n127 129.202
R638 vss.n129 vss.n128 129.202
R639 vss.n141 vss.n140 129.202
R640 vss.n140 vss.n139 129.202
R641 vss.n139 vss.n97 129.202
R642 vss.n333 vss.n97 129.202
R643 vss.n333 vss.n332 129.202
R644 vss.n330 vss.n96 124.832
R645 vss.n331 vss.n99 124.675
R646 vss.n317 vss.n104 122.373
R647 vss.n257 vss.n99 116.883
R648 vss.n261 vss.n257 116.883
R649 vss.n264 vss.n262 116.883
R650 vss.n264 vss.n263 116.883
R651 vss.n234 vss.n233 116.883
R652 vss.n244 vss.n234 116.883
R653 vss.n243 vss.n242 116.883
R654 vss.n242 vss.n235 116.883
R655 vss.n362 vss.n49 94.0779
R656 vss.n364 vss.n46 93.8579
R657 vss.n362 vss.t44 92.1964
R658 vss.n279 vss.t64 90.1798
R659 vss.n17 vss.n16 89.9525
R660 vss.n129 vss.t63 87.5698
R661 vss.t32 vss.n261 76.6239
R662 vss.n351 vss.n54 76.3222
R663 vss.n203 vss.n55 76.3222
R664 vss.n210 vss.n56 76.3222
R665 vss.n191 vss.n57 76.3222
R666 vss.n184 vss.n58 76.3222
R667 vss.n329 vss.n328 76.3222
R668 vss.n112 vss.n68 76.3222
R669 vss.n168 vss.n67 76.3222
R670 vss.n174 vss.n66 76.3222
R671 vss.n162 vss.n65 76.3222
R672 vss.n155 vss.n64 76.3222
R673 vss.n347 vss.n346 76.3222
R674 vss.n346 vss.n62 76.3222
R675 vss.n161 vss.n64 76.3222
R676 vss.n175 vss.n65 76.3222
R677 vss.n169 vss.n66 76.3222
R678 vss.n69 vss.n67 76.3222
R679 vss.n354 vss.n53 76.3222
R680 vss.n190 vss.n58 76.3222
R681 vss.n211 vss.n57 76.3222
R682 vss.n202 vss.n56 76.3222
R683 vss.n197 vss.n55 76.3222
R684 vss.n352 vss.n351 76.3222
R685 vss.n328 vss.n101 76.3222
R686 vss.n117 vss.n112 76.3222
R687 vss.n152 vss.n80 74.5978
R688 vss.n199 vss.n80 74.5978
R689 vss.n353 vss.t63 72.3318
R690 vss.t42 vss.n243 71.4291
R691 vss.n338 vss.n337 69.3109
R692 vss.n338 vss.n91 69.3109
R693 vss.n29 vss.n26 68.9197
R694 vss.n293 vss.n31 68.8547
R695 vss.n30 vss.n29 67.4522
R696 vss.n378 vss.n26 67.2825
R697 vss.n281 vss.n22 66.5677
R698 vss.t68 vss.n79 65.8183
R699 vss.t68 vss.n77 65.8183
R700 vss.t68 vss.n75 65.8183
R701 vss.t68 vss.n82 65.8183
R702 vss.t68 vss.n83 65.8183
R703 vss.t68 vss.n84 65.8183
R704 vss.t68 vss.n85 65.8183
R705 vss.t68 vss.n78 65.8183
R706 vss.t68 vss.n76 65.8183
R707 vss.t68 vss.n74 65.8183
R708 vss.n339 vss.t68 65.8183
R709 vss.t68 vss.n87 65.8183
R710 vss.t68 vss.n88 65.8183
R711 vss.t68 vss.n89 65.8183
R712 vss.t68 vss.n90 65.8183
R713 vss.n48 vss.n46 65.0005
R714 vss.n281 vss.n48 65.0005
R715 vss.n359 vss.n47 65.0005
R716 vss.n278 vss.n47 65.0005
R717 vss.n263 vss.t63 61.0395
R718 vss.t68 vss.n338 57.8461
R719 vss.n355 vss.n52 56.3995
R720 vss.n40 vss.n39 56.2007
R721 vss.n233 vss.t63 55.8447
R722 vss.t68 vss.n80 55.2026
R723 vss.n299 vss.n296 55.1712
R724 vss.n41 vss.n38 54.0035
R725 vss.n298 vss.n297 53.9338
R726 vss.n87 vss.n72 53.3664
R727 vss.n123 vss.n88 53.3664
R728 vss.n145 vss.n89 53.3664
R729 vss.n134 vss.n90 53.3664
R730 vss.n340 vss.n339 53.3664
R731 vss.n171 vss.n74 53.3664
R732 vss.n165 vss.n76 53.3664
R733 vss.n158 vss.n78 53.3664
R734 vss.n206 vss.n85 53.3664
R735 vss.n193 vss.n84 53.3664
R736 vss.n186 vss.n83 53.3664
R737 vss.n182 vss.n82 53.3664
R738 vss.n267 vss.n75 53.3664
R739 vss.n253 vss.n77 53.3664
R740 vss.n248 vss.n79 53.3664
R741 vss.n229 vss.n79 53.3664
R742 vss.n249 vss.n77 53.3664
R743 vss.n252 vss.n75 53.3664
R744 vss.n187 vss.n82 53.3664
R745 vss.n194 vss.n83 53.3664
R746 vss.n207 vss.n84 53.3664
R747 vss.n200 vss.n85 53.3664
R748 vss.n153 vss.n78 53.3664
R749 vss.n157 vss.n76 53.3664
R750 vss.n164 vss.n74 53.3664
R751 vss.n339 vss.n73 53.3664
R752 vss.n122 vss.n87 53.3664
R753 vss.n146 vss.n88 53.3664
R754 vss.n133 vss.n89 53.3664
R755 vss.n92 vss.n90 53.3664
R756 vss.n4 vss.n1 53.1823
R757 vss.t13 vss.n4 53.1823
R758 vss.n3 vss.n2 53.1823
R759 vss.t13 vss.n3 53.1823
R760 vss.n219 vss.n45 52.0418
R761 vss.n378 vss.n377 51.5266
R762 vss.n244 vss.t42 45.455
R763 vss.n385 vss.n384 42.0571
R764 vss.n141 vss.t63 41.6318
R765 vss.n8 vss.n2 41.1681
R766 vss.n262 vss.t32 40.2602
R767 vss.n305 vss.n35 39.7638
R768 vss.n303 vss.n287 39.511
R769 vss.n376 vss.n31 37.2591
R770 vss.n358 vss.n45 36.755
R771 vss.n377 vss.n376 36.6884
R772 vss.n29 vss.n28 36.563
R773 vss.n379 vss.n378 36.563
R774 vss.n314 vss.n312 35.7499
R775 vss.n384 vss.n383 34.4123
R776 vss.n383 vss.n382 34.4123
R777 vss.n15 vss.n14 34.4123
R778 vss.n14 vss.n13 34.4123
R779 vss.n293 vss.n292 32.5005
R780 vss.n306 vss.n305 32.5005
R781 vss.n307 vss.n306 32.5005
R782 vss.n325 vss.n324 32.1396
R783 vss.n1 vss.t14 30.8834
R784 vss.n283 vss.t15 30.0026
R785 vss.n235 vss.t36 29.8706
R786 vss.t34 vss.t78 29.1645
R787 vss.t54 vss.t75 29.1645
R788 vss.t58 vss.t77 29.1645
R789 vss.t38 vss.t76 29.1645
R790 vss.t52 vss.t9 29.1645
R791 vss.t59 vss.t8 29.1645
R792 vss.t48 vss.t6 29.1645
R793 vss.t40 vss.t5 29.1645
R794 vss.t61 vss.t7 29.1645
R795 vss.t17 vss.t44 29.1645
R796 vss.t16 vss.t56 29.1645
R797 vss.t19 vss.t65 29.1645
R798 vss.t15 vss.t50 29.0651
R799 vss.t62 vss.t24 29.0651
R800 vss.t26 vss.t22 29.0651
R801 vss.n312 vss.t76 27.2829
R802 vss.t7 vss.n49 27.2829
R803 vss.n218 vss.t27 26.5035
R804 vss.n357 vss.n356 25.5303
R805 vss.n271 vss.t33 25.0376
R806 vss.n359 vss.n358 23.4151
R807 vss.n18 vss.n17 23.0405
R808 vss.n27 vss.t20 22.4758
R809 vss.n218 vss.n217 20.6876
R810 vss.n221 vss.n216 20.6876
R811 vss.n222 vss.n215 20.6876
R812 vss.n320 vss.n272 20.6683
R813 vss.n319 vss.n273 20.6683
R814 vss.n275 vss.n274 20.6683
R815 vss.n44 vss.n43 20.6683
R816 vss.n16 vss.n15 18.7337
R817 vss.n15 vss.n9 16.3845
R818 vss.n373 vss.n34 15.5385
R819 vss.n282 vss.t21 15.0016
R820 vss.n277 vss.n276 14.6255
R821 vss.n282 vss.n277 14.6255
R822 vss.n325 vss.n98 14.6255
R823 vss.n331 vss.n98 14.6255
R824 vss.t64 vss.t74 14.5716
R825 vss.t18 vss.t30 14.5576
R826 vss.n377 vss.n30 14.2889
R827 vss.n11 vss.n9 11.9393
R828 vss.n12 vss.n11 11.9393
R829 vss.n20 vss.n19 11.9393
R830 vss.n21 vss.n20 11.9393
R831 vss.n296 vss.t11 11.6005
R832 vss.n296 vss.t67 11.6005
R833 vss.n297 vss.t2 11.6005
R834 vss.n297 vss.t73 11.6005
R835 vss.n38 vss.t3 11.6005
R836 vss.n38 vss.t72 11.6005
R837 vss.n39 vss.t79 11.6005
R838 vss.n39 vss.t70 11.6005
R839 vss.n295 vss.n294 10.5495
R840 vss.n16 vss.n1 10.0532
R841 vss.n345 vss.n63 9.36638
R842 vss.n375 vss.n32 9.35616
R843 vss.n301 vss.n287 9.3005
R844 vss.n372 vss.n371 9.3005
R845 vss.n286 vss.n36 9.3005
R846 vss.n291 vss.t10 8.47308
R847 vss.n18 vss.n6 7.5005
R848 vss.n10 vss.n6 7.5005
R849 vss.n7 vss.n5 7.5005
R850 vss.n10 vss.n5 7.5005
R851 vss.n364 vss.n363 7.313
R852 vss.n363 vss.n362 7.313
R853 vss.n361 vss.n360 7.313
R854 vss.n362 vss.n361 7.313
R855 vss.n324 vss.n323 6.9005
R856 vss.n322 vss.n104 6.9005
R857 vss.t46 vss.n278 6.57608
R858 vss.n365 vss.n45 6.51916
R859 vss.n316 vss.n315 6.15839
R860 vss.n315 vss.n314 6.15839
R861 vss.n313 vss.n50 6.15839
R862 vss.n314 vss.n313 6.15839
R863 vss.n343 vss.n342 4.90263
R864 vss.n349 vss.n348 4.90263
R865 vss.n121 vss.n120 4.88977
R866 vss.n125 vss.n124 4.88977
R867 vss.n143 vss.n108 4.88977
R868 vss.n135 vss.n132 4.88977
R869 vss.n137 vss.n136 4.88977
R870 vss.n336 vss.n93 4.88977
R871 vss.n294 vss.n285 4.8755
R872 vss.n290 vss.n285 4.8755
R873 vss.n284 vss.n34 4.8755
R874 vss.n290 vss.n284 4.8755
R875 vss.n335 vss.n94 4.65477
R876 vss.n100 vss.n94 4.57193
R877 vss.n301 vss.n289 4.5005
R878 vss.n371 vss.n370 4.5005
R879 vss.n369 vss.n36 4.5005
R880 vss.n272 vss.t43 4.3505
R881 vss.n272 vss.t37 4.3505
R882 vss.n273 vss.t35 4.3505
R883 vss.n273 vss.t55 4.3505
R884 vss.n274 vss.t49 4.3505
R885 vss.n274 vss.t41 4.3505
R886 vss.n43 vss.t31 4.3505
R887 vss.n43 vss.t51 4.3505
R888 vss.n217 vss.t45 4.3505
R889 vss.n217 vss.t57 4.3505
R890 vss.n216 vss.t39 4.3505
R891 vss.n216 vss.t53 4.3505
R892 vss.n215 vss.t29 4.3505
R893 vss.n215 vss.t47 4.3505
R894 vss.n119 vss.n70 4.23054
R895 vss.n375 vss.n374 4.1842
R896 vss.n37 vss.n33 4.11666
R897 vss.n323 vss.n271 4.10351
R898 vss.n327 vss.n326 3.9624
R899 vss.n201 vss.n198 3.81327
R900 vss.n205 vss.n204 3.81327
R901 vss.n208 vss.n196 3.81327
R902 vss.n209 vss.n179 3.81327
R903 vss.n212 vss.n195 3.81327
R904 vss.n192 vss.n180 3.81327
R905 vss.n189 vss.n188 3.81327
R906 vss.n185 vss.n183 3.81327
R907 vss.n372 vss.n35 3.76521
R908 vss.n385 vss.n1 3.71562
R909 vss.n111 vss.n70 3.70433
R910 vss.n219 vss.n50 3.60613
R911 vss.n148 vss.n147 3.51638
R912 vss.n107 vss.n106 3.35157
R913 vss.n386 vss.n0 3.33015
R914 vss.n368 vss.n0 3.1874
R915 vss.n350 vss.n60 3.15965
R916 vss.n341 vss.n71 2.7239
R917 vss.n170 vss.n167 2.7239
R918 vss.n173 vss.n172 2.7239
R919 vss.n166 vss.n163 2.7239
R920 vss.n160 vss.n150 2.7239
R921 vss.n159 vss.n156 2.7239
R922 vss.n154 vss.n151 2.7239
R923 vss.n348 vss.n61 2.7239
R924 vss.n367 vss.n366 2.49883
R925 vss.n301 vss.n300 2.34663
R926 vss.n323 vss.n322 2.28754
R927 vss.n367 vss.n44 2.27913
R928 vss.n342 vss.n341 2.17922
R929 vss.n167 vss.n71 2.17922
R930 vss.n172 vss.n170 2.17922
R931 vss.n173 vss.n149 2.17922
R932 vss.n176 vss.n166 2.17922
R933 vss.n163 vss.n150 2.17922
R934 vss.n160 vss.n159 2.17922
R935 vss.n156 vss.n154 2.17922
R936 vss.n151 vss.n61 2.17922
R937 vss.n240 vss.n239 2.17819
R938 vss.n370 vss.n41 2.11938
R939 vss.n270 vss.n269 1.89157
R940 vss.n350 vss.n349 1.85241
R941 vss.n259 vss.n258 1.79105
R942 vss.n266 vss.n225 1.79105
R943 vss.n255 vss.n254 1.79105
R944 vss.n247 vss.n228 1.79105
R945 vss.n246 vss.n230 1.79105
R946 vss.n238 vss.n237 1.79105
R947 vss vss.n250 1.76685
R948 vss.n41 vss.n40 1.74237
R949 vss.n386 vss.n385 1.7255
R950 vss.n366 vss 1.6569
R951 vss.n177 vss.n176 1.63454
R952 vss.n356 vss.n51 1.62167
R953 vss.n144 vss.n107 1.5387
R954 vss.n343 vss.n70 1.52561
R955 vss.n178 vss.n148 1.51978
R956 vss.n222 vss.n221 1.46641
R957 vss.n220 vss.n218 1.43895
R958 vss.n326 vss.n103 1.37971
R959 vss.n148 vss.n105 1.37389
R960 vss.n304 vss.n303 1.30961
R961 vss.n298 vss.n289 1.21619
R962 vss.n269 vss.n224 1.21033
R963 vss.n327 vss.n102 1.11796
R964 vss.n198 vss.n60 1.08986
R965 vss.n204 vss.n201 1.08986
R966 vss.n205 vss.n196 1.08986
R967 vss.n209 vss.n208 1.08986
R968 vss.n195 vss.n192 1.08986
R969 vss.n189 vss.n180 1.08986
R970 vss.n188 vss.n185 1.08986
R971 vss.n183 vss.n181 1.08986
R972 vss.n181 vss.n51 1.08986
R973 vss.n177 vss.n149 1.08986
R974 vss.n305 vss.n304 1.06085
R975 vss.n275 vss.n44 0.998567
R976 vss.n320 vss.n319 0.997923
R977 vss.n299 vss.n298 0.995892
R978 vss.n376 vss.n375 0.874635
R979 vss.n213 vss.n179 0.871989
R980 vss.n239 vss.n51 0.823184
R981 vss.n214 vss.n178 0.764974
R982 vss.n286 vss.n35 0.684992
R983 vss.n223 vss.n214 0.653909
R984 vss.n321 vss.n320 0.633876
R985 vss.n178 vss.n177 0.596304
R986 vss.n214 vss.n213 0.59175
R987 vss.n269 vss.n268 0.581218
R988 vss.t36 vss.t63 0.545594
R989 vss.n223 vss.n222 0.539326
R990 vss.n317 vss.n316 0.532356
R991 vss.n318 vss.n275 0.528206
R992 vss.n288 vss.n42 0.497949
R993 vss.n302 vss.n37 0.484781
R994 vss.n319 vss.n318 0.469572
R995 vss.n270 vss.n223 0.452516
R996 vss.n302 vss.n301 0.446546
R997 vss.n368 vss.n367 0.40709
R998 vss.n369 vss.n368 0.389161
R999 vss.n259 vss.n103 0.387646
R1000 vss.n258 vss.n224 0.387646
R1001 vss.n268 vss.n266 0.387646
R1002 vss.n255 vss.n225 0.387646
R1003 vss.n250 vss.n228 0.387646
R1004 vss.n247 vss.n246 0.387646
R1005 vss.n237 vss.n230 0.387646
R1006 vss.n240 vss.n238 0.387646
R1007 vss.t12 vss.t69 0.36604
R1008 vss.t4 vss.t0 0.36604
R1009 vss.n322 vss.n321 0.343093
R1010 vss.n303 vss.n302 0.32741
R1011 vss.n254 vss 0.266663
R1012 vss.n365 vss.n364 0.222008
R1013 vss.n213 vss.n212 0.218372
R1014 vss.n32 vss.n31 0.205848
R1015 vss.n369 vss.n42 0.141656
R1016 vss.n17 vss.n0 0.139042
R1017 vss.n302 vss.n42 0.1255
R1018 vss vss.n251 0.121483
R1019 vss vss.n386 0.120187
R1020 vss.n220 vss.n219 0.0987955
R1021 vss.n271 vss.n270 0.0952653
R1022 vss.n374 vss.n373 0.0850455
R1023 vss.n321 vss 0.0849072
R1024 vss.n288 vss 0.0796284
R1025 vss.n318 vss.n317 0.0736577
R1026 vss.n366 vss.n365 0.0596905
R1027 vss.n120 vss.n119 0.0554356
R1028 vss.n125 vss.n121 0.0554356
R1029 vss.n124 vss.n105 0.0554356
R1030 vss.n147 vss.n106 0.0554356
R1031 vss.n144 vss.n143 0.0554356
R1032 vss.n132 vss.n108 0.0554356
R1033 vss.n137 vss.n135 0.0554356
R1034 vss.n136 vss.n93 0.0554356
R1035 vss.n336 vss.n335 0.0554356
R1036 vss.n102 vss.n100 0.0512937
R1037 vss.n371 vss.n37 0.0386737
R1038 vss.n40 vss.n33 0.0370854
R1039 vss.n374 vss.n33 0.0287609
R1040 vss.n300 vss.n295 0.0286818
R1041 vss.n221 vss.n220 0.0279621
R1042 vss.n289 vss.n288 0.0274495
R1043 vss.n251 vss 0.0246966
R1044 vss.n370 vss.n369 0.0152996
R1045 vss.n300 vss.n299 0.0126951
R1046 vss.n371 vss.n36 0.00424252
R1047 OTA_vref_0.OTA_vref_stage2_0.vr.n0 OTA_vref_0.OTA_vref_stage2_0.vr.t3 651.943
R1048 OTA_vref_0.OTA_vref_stage2_0.vr.n18 OTA_vref_0.OTA_vref_stage2_0.vr.t1 651.678
R1049 OTA_vref_0.OTA_vref_stage2_0.vr.n20 OTA_vref_0.OTA_vref_stage2_0.vr.t22 60.1752
R1050 OTA_vref_0.OTA_vref_stage2_0.vr.n19 OTA_vref_0.OTA_vref_stage2_0.vr.t25 60.1752
R1051 OTA_vref_0.OTA_vref_stage2_0.vr.n4 OTA_vref_0.OTA_vref_stage2_0.vr.t8 28.5589
R1052 OTA_vref_0.OTA_vref_stage2_0.vr.n7 OTA_vref_0.OTA_vref_stage2_0.vr.t10 27.6016
R1053 OTA_vref_0.OTA_vref_stage2_0.vr.n21 OTA_vref_0.OTA_vref_stage2_0.vr.t21 26.8562
R1054 OTA_vref_0.OTA_vref_stage2_0.vr.n21 OTA_vref_0.OTA_vref_stage2_0.vr.t23 26.0492
R1055 OTA_vref_0.OTA_vref_stage2_0.vr.n22 OTA_vref_0.OTA_vref_stage2_0.vr.t20 26.0492
R1056 OTA_vref_0.OTA_vref_stage2_0.vr.n23 OTA_vref_0.OTA_vref_stage2_0.vr.t26 26.0492
R1057 OTA_vref_0.OTA_vref_stage2_0.vr.n24 OTA_vref_0.OTA_vref_stage2_0.vr.t24 26.0492
R1058 OTA_vref_0.OTA_vref_stage2_0.vr.n11 OTA_vref_0.OTA_vref_stage2_0.vr.n10 24.2089
R1059 OTA_vref_0.OTA_vref_stage2_0.vr.n12 OTA_vref_0.OTA_vref_stage2_0.vr.n8 23.2516
R1060 OTA_vref_0.OTA_vref_stage2_0.vr.n11 OTA_vref_0.OTA_vref_stage2_0.vr.n9 23.2516
R1061 OTA_vref_0.OTA_vref_stage2_0.vr.n6 OTA_vref_0.OTA_vref_stage2_0.vr.n1 23.2516
R1062 OTA_vref_0.OTA_vref_stage2_0.vr.n5 OTA_vref_0.OTA_vref_stage2_0.vr.n2 23.2516
R1063 OTA_vref_0.OTA_vref_stage2_0.vr.n4 OTA_vref_0.OTA_vref_stage2_0.vr.n3 23.2516
R1064 OTA_vref_0.OTA_vref_stage2_0.vr.n14 OTA_vref_0.OTA_vref_stage2_0.vr.n13 23.2516
R1065 OTA_vref_0.OTA_vref_stage2_0.vr.n17 OTA_vref_0.OTA_vref_stage2_0.vr.t0 23
R1066 OTA_vref_0.OTA_vref_stage2_0.vr.n0 OTA_vref_0.OTA_vref_stage2_0.vr.t2 23
R1067 OTA_vref_0.OTA_vref_stage2_0.vr.n8 OTA_vref_0.OTA_vref_stage2_0.vr.t15 4.3505
R1068 OTA_vref_0.OTA_vref_stage2_0.vr.n8 OTA_vref_0.OTA_vref_stage2_0.vr.t7 4.3505
R1069 OTA_vref_0.OTA_vref_stage2_0.vr.n9 OTA_vref_0.OTA_vref_stage2_0.vr.t4 4.3505
R1070 OTA_vref_0.OTA_vref_stage2_0.vr.n9 OTA_vref_0.OTA_vref_stage2_0.vr.t18 4.3505
R1071 OTA_vref_0.OTA_vref_stage2_0.vr.n10 OTA_vref_0.OTA_vref_stage2_0.vr.t12 4.3505
R1072 OTA_vref_0.OTA_vref_stage2_0.vr.n10 OTA_vref_0.OTA_vref_stage2_0.vr.t5 4.3505
R1073 OTA_vref_0.OTA_vref_stage2_0.vr.n1 OTA_vref_0.OTA_vref_stage2_0.vr.t9 4.3505
R1074 OTA_vref_0.OTA_vref_stage2_0.vr.n1 OTA_vref_0.OTA_vref_stage2_0.vr.t14 4.3505
R1075 OTA_vref_0.OTA_vref_stage2_0.vr.n2 OTA_vref_0.OTA_vref_stage2_0.vr.t11 4.3505
R1076 OTA_vref_0.OTA_vref_stage2_0.vr.n2 OTA_vref_0.OTA_vref_stage2_0.vr.t16 4.3505
R1077 OTA_vref_0.OTA_vref_stage2_0.vr.n3 OTA_vref_0.OTA_vref_stage2_0.vr.t13 4.3505
R1078 OTA_vref_0.OTA_vref_stage2_0.vr.n3 OTA_vref_0.OTA_vref_stage2_0.vr.t6 4.3505
R1079 OTA_vref_0.OTA_vref_stage2_0.vr.n13 OTA_vref_0.OTA_vref_stage2_0.vr.t19 4.3505
R1080 OTA_vref_0.OTA_vref_stage2_0.vr.n13 OTA_vref_0.OTA_vref_stage2_0.vr.t17 4.3505
R1081 OTA_vref_0.OTA_vref_stage2_0.vr.n16 OTA_vref_0.OTA_vref_stage2_0.vr.n15 3.8934
R1082 OTA_vref_0.OTA_vref_stage2_0.vr.n22 OTA_vref_0.OTA_vref_stage2_0.vr.n21 2.80213
R1083 OTA_vref_0.OTA_vref_stage2_0.vr.n24 OTA_vref_0.OTA_vref_stage2_0.vr.n23 2.76952
R1084 OTA_vref_0.OTA_vref_stage2_0.vr.n23 OTA_vref_0.OTA_vref_stage2_0.vr.n22 2.72333
R1085 OTA_vref_0.OTA_vref_stage2_0.vr.n15 OTA_vref_0.OTA_vref_stage2_0.vr.n14 1.06728
R1086 OTA_vref_0.OTA_vref_stage2_0.vr.n7 OTA_vref_0.OTA_vref_stage2_0.vr.n6 0.957816
R1087 OTA_vref_0.OTA_vref_stage2_0.vr.n6 OTA_vref_0.OTA_vref_stage2_0.vr.n5 0.957816
R1088 OTA_vref_0.OTA_vref_stage2_0.vr.n5 OTA_vref_0.OTA_vref_stage2_0.vr.n4 0.957816
R1089 OTA_vref_0.OTA_vref_stage2_0.vr.n14 OTA_vref_0.OTA_vref_stage2_0.vr.n12 0.957816
R1090 OTA_vref_0.OTA_vref_stage2_0.vr.n12 OTA_vref_0.OTA_vref_stage2_0.vr.n11 0.957816
R1091 OTA_vref_0.OTA_vref_stage2_0.vr.n19 OTA_vref_0.OTA_vref_stage2_0.vr.n18 0.774957
R1092 OTA_vref_0.OTA_vref_stage2_0.vr OTA_vref_0.OTA_vref_stage2_0.vr.n20 0.660826
R1093 OTA_vref_0.OTA_vref_stage2_0.vr OTA_vref_0.OTA_vref_stage2_0.vr.n24 0.617348
R1094 OTA_vref_0.OTA_vref_stage2_0.vr.n15 OTA_vref_0.OTA_vref_stage2_0.vr.n7 0.577487
R1095 OTA_vref_0.OTA_vref_stage2_0.vr.n20 OTA_vref_0.OTA_vref_stage2_0.vr.n19 0.36463
R1096 OTA_vref_0.OTA_vref_stage2_0.vr.n18 OTA_vref_0.OTA_vref_stage2_0.vr.n17 0.269439
R1097 OTA_vref_0.OTA_vref_stage2_0.vr.n17 OTA_vref_0.OTA_vref_stage2_0.vr.n16 0.240192
R1098 OTA_vref_0.OTA_vref_stage2_0.vr.n16 OTA_vref_0.OTA_vref_stage2_0.vr.n0 0.216951
R1099 vin_p.n0 vin_p.t0 21.6012
R1100 vin_p.n0 vin_p.t1 8.85318
R1101 vin_p vin_p.n0 2.55816
R1102 OTA_stage2_0.vd2.t0 OTA_stage2_0.vd2.t2 134.761
R1103 OTA_stage2_0.vd2.t0 OTA_stage2_0.vd2.t1 134.73
R1104 OTA_stage2_0.vd2.t0 OTA_stage2_0.vd2.t6 129.905
R1105 OTA_stage2_0.vd2.t0 OTA_stage2_0.vd2.t4 122.688
R1106 OTA_stage2_0.vd2.t0 OTA_stage2_0.vd2.t3 122.213
R1107 OTA_stage2_0.vd2.t0 OTA_stage2_0.vd2.t5 122.213
R1108 OTA_vref_0.vb1.n1 OTA_vref_0.vb1.n2 71.7516
R1109 OTA_vref_0.vb1.n1 OTA_vref_0.vb1.n3 70.9453
R1110 OTA_vref_0.vb1.n1 OTA_vref_0.vb1.n4 70.9453
R1111 OTA_vref_0.vb1.n0 OTA_vref_0.vb1.t7 68.1062
R1112 OTA_vref_0.vb1.n0 OTA_vref_0.vb1.t6 67.5138
R1113 OTA_vref_0.vb1.n0 OTA_vref_0.vb1.t9 67.5138
R1114 OTA_vref_0.vb1.n0 OTA_vref_0.vb1.t8 67.5138
R1115 OTA_vref_0.vb1.n2 OTA_vref_0.vb1.t2 17.4005
R1116 OTA_vref_0.vb1.n2 OTA_vref_0.vb1.t5 17.4005
R1117 OTA_vref_0.vb1.n3 OTA_vref_0.vb1.t1 17.4005
R1118 OTA_vref_0.vb1.n3 OTA_vref_0.vb1.t0 17.4005
R1119 OTA_vref_0.vb1.n4 OTA_vref_0.vb1.t4 17.4005
R1120 OTA_vref_0.vb1.n4 OTA_vref_0.vb1.t3 17.4005
R1121 OTA_stage2_0.vb1 OTA_vref_0.vb1.n0 10.0221
R1122 OTA_vref_0.OTA_vref_stage2_0.vb1 OTA_vref_0.vb1.n1 8.73695
R1123 OTA_vref_0.OTA_vref_stage2_0.vb1 OTA_stage2_0.vb1 6.72684
R1124 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t3 138.714
R1125 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t4 136.073
R1126 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t7 122.216
R1127 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t5 122.216
R1128 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t6 121.828
R1129 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t8 121.828
R1130 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t0 19.5045
R1131 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t1 17.559
R1132 OTA_stage2_0.vd1.n0 OTA_stage2_0.vd1.t2 16.4891
R1133 vo.n3 vo.t7 72.7606
R1134 vo.n4 vo.t8 71.6732
R1135 vo.n7 vo.n6 62.1978
R1136 vo.n5 vo.t5 52.9855
R1137 vo.n0 vo.t3 19.4751
R1138 vo.n0 vo.t2 18.6511
R1139 vo.n2 vo.n1 15.6099
R1140 vo.n6 vo.t6 11.6005
R1141 vo.n6 vo.t0 11.6005
R1142 vo.n4 vo.n3 2.48505
R1143 vo.n1 vo.t1 1.90483
R1144 vo.n1 vo.t4 1.90483
R1145 vo.n2 vo.n0 1.32214
R1146 vo.n3 vo.n2 1.28407
R1147 vo.n7 vo.n5 0.307843
R1148 vo vo.n7 0.0135556
R1149 vo.n5 vo.n4 0.00787255
R1150 a_959_2177.n4 a_959_2177.t11 36.4777
R1151 a_959_2177.n5 a_959_2177.t8 35.4327
R1152 a_959_2177.n4 a_959_2177.n3 31.3519
R1153 a_959_2177.n8 a_959_2177.n7 18.3035
R1154 a_959_2177.n2 a_959_2177.n1 18.303
R1155 a_959_2177.n9 a_959_2177.n8 17.2098
R1156 a_959_2177.n2 a_959_2177.n0 17.208
R1157 a_959_2177.n6 a_959_2177.n2 8.938
R1158 a_959_2177.n3 a_959_2177.t9 4.08121
R1159 a_959_2177.n3 a_959_2177.t10 4.08121
R1160 a_959_2177.n8 a_959_2177.n6 3.05142
R1161 a_959_2177.n6 a_959_2177.n5 2.2455
R1162 a_959_2177.n1 a_959_2177.t6 1.90483
R1163 a_959_2177.n1 a_959_2177.t2 1.90483
R1164 a_959_2177.n0 a_959_2177.t0 1.90483
R1165 a_959_2177.n0 a_959_2177.t5 1.90483
R1166 a_959_2177.n7 a_959_2177.t1 1.90483
R1167 a_959_2177.n7 a_959_2177.t7 1.90483
R1168 a_959_2177.n9 a_959_2177.t4 1.90483
R1169 a_959_2177.t3 a_959_2177.n9 1.90483
R1170 a_959_2177.n5 a_959_2177.n4 1.0455
R1171 vcc.n146 vcc.n19 17565.9
R1172 vcc.n148 vcc.n19 17565.9
R1173 vcc.n148 vcc.n20 17562.4
R1174 vcc.n146 vcc.n20 17562.4
R1175 vcc.n8 vcc.n5 16027.1
R1176 vcc.n10 vcc.n5 16027.1
R1177 vcc.n8 vcc.n6 16027.1
R1178 vcc.n10 vcc.n6 16027.1
R1179 vcc.n137 vcc.n121 6349.41
R1180 vcc.n137 vcc.n122 6349.41
R1181 vcc.n135 vcc.n121 6349.41
R1182 vcc.n135 vcc.n122 6349.41
R1183 vcc.n51 vcc.n45 3045.88
R1184 vcc.n51 vcc.n46 3045.88
R1185 vcc.n49 vcc.n45 3045.88
R1186 vcc.n49 vcc.n46 3045.88
R1187 vcc.n80 vcc.n79 2706.92
R1188 vcc.n95 vcc.n79 2701.93
R1189 vcc.n93 vcc.n92 2375
R1190 vcc.n92 vcc.n80 2327.31
R1191 vcc.n75 vcc.n32 2089.41
R1192 vcc.n72 vcc.n33 2089.41
R1193 vcc.n64 vcc.n37 2089.41
R1194 vcc.n67 vcc.n66 2089.41
R1195 vcc.n57 vcc.n41 2089.41
R1196 vcc.n60 vcc.n59 2089.41
R1197 vcc.n10 vcc.t25 1353.8
R1198 vcc.t22 vcc.n8 1317.74
R1199 vcc.n9 vcc.t22 1196.03
R1200 vcc.t25 vcc.n9 1159.97
R1201 vcc.n90 vcc.t4 653.497
R1202 vcc.t0 vcc.n80 616.96
R1203 vcc.n84 vcc.n83 599.49
R1204 vcc.t14 vcc.n49 538
R1205 vcc.n54 vcc.n43 524.801
R1206 vcc.n51 vcc.t10 524.534
R1207 vcc.n91 vcc.t0 519.274
R1208 vcc.t10 vcc.n50 441.339
R1209 vcc.n50 vcc.t14 427.875
R1210 vcc.n73 vcc.n32 426.346
R1211 vcc.n74 vcc.n33 426.346
R1212 vcc.n65 vcc.n64 426.346
R1213 vcc.n67 vcc.n36 426.346
R1214 vcc.n58 vcc.n57 426.346
R1215 vcc.n60 vcc.n39 426.346
R1216 vcc.n7 vcc.n4 415.628
R1217 vcc.n11 vcc.n4 405.284
R1218 vcc.t4 vcc.t12 387.817
R1219 vcc.n88 vcc.n87 300.267
R1220 vcc.n95 vcc.n94 268.39
R1221 vcc.n89 vcc.n78 253.333
R1222 vcc.n89 vcc.n88 248.246
R1223 vcc.n104 vcc.t17 231.287
R1224 vcc.n103 vcc.t3 231.287
R1225 vcc.n102 vcc.t9 231.287
R1226 vcc.n24 vcc.t11 231.273
R1227 vcc.n108 vcc.t15 231.273
R1228 vcc.t28 vcc.t30 216.05
R1229 vcc.t34 vcc.t32 216.05
R1230 vcc.n145 vcc.n16 209.422
R1231 vcc.n101 vcc.n26 202.453
R1232 vcc.t6 vcc.n90 198.105
R1233 vcc.n7 vcc.n3 183.016
R1234 vcc.n12 vcc.n11 176.572
R1235 vcc.t30 vcc.n121 174.992
R1236 vcc.t32 vcc.n122 174.992
R1237 vcc.n91 vcc.t6 168.089
R1238 vcc.n150 vcc.n17 157.375
R1239 vcc.n48 vcc.n47 128.981
R1240 vcc.n2 vcc.n0 120.891
R1241 vcc.n2 vcc.n1 119.76
R1242 vcc.n96 vcc.n78 118.118
R1243 vcc.n117 vcc.n116 116.722
R1244 vcc.n149 vcc.n18 115.912
R1245 vcc.n150 vcc.n149 108.909
R1246 vcc.n136 vcc.t28 108.025
R1247 vcc.n136 vcc.t34 108.025
R1248 vcc.n47 vcc.n43 103.507
R1249 vcc.n71 vcc.n30 101.719
R1250 vcc.n112 vcc.n111 87.9664
R1251 vcc.n112 vcc.n18 87.7954
R1252 vcc.n71 vcc.n70 82.4041
R1253 vcc.n62 vcc.n34 73.7015
R1254 vcc.n69 vcc.n34 72.4513
R1255 vcc.n125 vcc.n124 71.8902
R1256 vcc.t18 vcc.n146 71.3347
R1257 vcc.n134 vcc.n123 70.7824
R1258 vcc.n141 vcc.n21 65.6211
R1259 vcc.n40 vcc.n38 64.6513
R1260 vcc.n55 vcc.n40 64.1322
R1261 vcc.n88 vcc.n80 61.6672
R1262 vcc.n148 vcc.t20 60.8049
R1263 vcc.n97 vcc.n96 58.2536
R1264 vcc.n83 vcc.t1 57.1305
R1265 vcc.n83 vcc.t7 57.1305
R1266 vcc.n145 vcc.n144 55.3321
R1267 vcc.t21 vcc.t18 53.6285
R1268 vcc.t20 vcc.t19 53.6285
R1269 vcc.n138 vcc.n120 50.9389
R1270 vcc.n93 vcc.n78 46.2505
R1271 vcc.n53 vcc.n44 45.9062
R1272 vcc.n48 vcc.n44 45.8838
R1273 vcc.n53 vcc.n52 38.0921
R1274 vcc.n77 vcc.n30 36.2672
R1275 vcc.n52 vcc.n43 35.1619
R1276 vcc.n94 vcc.n93 33.6365
R1277 vcc.n128 vcc.n126 32.1789
R1278 vcc.t19 vcc.n147 32.0794
R1279 vcc.n128 vcc.n127 32.0774
R1280 vcc.n49 vcc.n48 30.8799
R1281 vcc.n52 vcc.n51 30.8338
R1282 vcc.n57 vcc.n56 30.8338
R1283 vcc.n64 vcc.n63 30.8338
R1284 vcc.n61 vcc.n60 30.8338
R1285 vcc.n32 vcc.n31 30.8338
R1286 vcc.n68 vcc.n67 30.8338
R1287 vcc.n33 vcc.n30 30.8338
R1288 vcc.n96 vcc.n95 30.8338
R1289 vcc.n94 vcc.t12 30.7518
R1290 vcc.n117 vcc.n21 30.7043
R1291 vcc.n139 vcc.n138 30.0503
R1292 vcc.n139 vcc.n119 29.6052
R1293 vcc.n26 vcc.t5 28.5655
R1294 vcc.n26 vcc.t13 28.5655
R1295 vcc.n76 vcc.n75 23.1255
R1296 vcc.n37 vcc.n35 23.1255
R1297 vcc.n42 vcc.n41 23.1255
R1298 vcc.n59 vcc.n40 23.1255
R1299 vcc.n66 vcc.n34 23.1255
R1300 vcc.n72 vcc.n71 23.1255
R1301 vcc.n147 vcc.t21 21.5497
R1302 vcc.n75 vcc.n74 18.2059
R1303 vcc.n37 vcc.n36 18.2059
R1304 vcc.n41 vcc.n39 18.2059
R1305 vcc.n59 vcc.n58 18.2059
R1306 vcc.n66 vcc.n65 18.2059
R1307 vcc.n73 vcc.n72 18.2059
R1308 vcc.n1 vcc.t24 15.8699
R1309 vcc.n1 vcc.t27 15.8699
R1310 vcc.n0 vcc.t23 15.8699
R1311 vcc.n0 vcc.t26 15.8699
R1312 vcc.n98 vcc.n97 13.5977
R1313 vcc.n81 vcc.n29 12.7275
R1314 vcc.n97 vcc.n77 12.0301
R1315 vcc.n92 vcc.n89 11.563
R1316 vcc.n92 vcc.n91 11.563
R1317 vcc.n47 vcc.n46 10.8829
R1318 vcc.n50 vcc.n46 10.8829
R1319 vcc.n45 vcc.n44 10.8829
R1320 vcc.n50 vcc.n45 10.8829
R1321 vcc.n77 vcc.n76 10.3636
R1322 vcc.n11 vcc.n10 10.2783
R1323 vcc.n8 vcc.n7 10.2783
R1324 vcc.n63 vcc.n35 9.97982
R1325 vcc.n70 vcc.n69 9.87337
R1326 vcc.n76 vcc.n31 9.86377
R1327 vcc.n68 vcc.n35 9.83647
R1328 vcc.n56 vcc.n42 9.75729
R1329 vcc.n84 vcc 9.63246
R1330 vcc.n62 vcc.n61 9.62493
R1331 vcc.n42 vcc.n25 9.57855
R1332 vcc.n116 vcc.n115 9.34567
R1333 vcc.n99 vcc.n98 9.3005
R1334 vcc.n29 vcc.n28 9.3005
R1335 vcc.n133 vcc.n132 9.3005
R1336 vcc.n142 vcc.n141 9.3005
R1337 vcc.n113 vcc.n112 9.3005
R1338 vcc.n55 vcc.n54 9.07124
R1339 vcc.n124 vcc.n122 8.04398
R1340 vcc.n123 vcc.n121 8.04398
R1341 vcc.n81 vcc.n79 7.4005
R1342 vcc.n90 vcc.n79 7.4005
R1343 vcc vcc.n101 7.20708
R1344 vcc.n135 vcc.n134 7.11588
R1345 vcc.n136 vcc.n135 7.11588
R1346 vcc.n138 vcc.n137 7.11588
R1347 vcc.n137 vcc.n136 7.11588
R1348 vcc.n144 vcc.n21 6.56253
R1349 vcc.n111 vcc.n20 5.44168
R1350 vcc.n147 vcc.n20 5.44168
R1351 vcc.n19 vcc.n17 5.44168
R1352 vcc.n147 vcc.n19 5.44168
R1353 vcc.n134 vcc.n133 4.82369
R1354 vcc.n74 vcc.t8 4.71965
R1355 vcc.t8 vcc.n73 4.71965
R1356 vcc.t2 vcc.n36 4.71965
R1357 vcc.n65 vcc.t2 4.71965
R1358 vcc.t16 vcc.n39 4.71965
R1359 vcc.n58 vcc.t16 4.71965
R1360 vcc.n114 vcc.n113 4.5005
R1361 vcc.n123 vcc.n120 4.48345
R1362 vcc.n116 vcc.n22 4.42232
R1363 vcc.n126 vcc.t31 4.08121
R1364 vcc.n126 vcc.t29 4.08121
R1365 vcc.n127 vcc.t35 4.08121
R1366 vcc.n127 vcc.t33 4.08121
R1367 vcc.n107 vcc.n106 3.76209
R1368 vcc.n100 vcc.n99 2.2505
R1369 vcc.n133 vcc.n125 1.94833
R1370 vcc.n111 vcc.n22 1.86232
R1371 vcc.n152 vcc.n151 1.85361
R1372 vcc.n108 vcc.n107 1.80651
R1373 vcc.n146 vcc.n145 1.66717
R1374 vcc.n149 vcc.n148 1.66717
R1375 vcc.n6 vcc.n4 1.63767
R1376 vcc.n9 vcc.n6 1.63767
R1377 vcc.n5 vcc.n3 1.63767
R1378 vcc.n9 vcc.n5 1.63767
R1379 vcc.n140 vcc.n139 1.6211
R1380 vcc.n15 vcc.n14 1.42554
R1381 vcc.n98 vcc.n29 1.27753
R1382 vcc.n13 vcc 1.27612
R1383 vcc.n154 vcc.n15 1.21717
R1384 vcc.n17 vcc.n16 1.20392
R1385 vcc.n14 vcc.n2 1.20189
R1386 vcc.n124 vcc.n119 1.19816
R1387 vcc.n113 vcc.n110 1.19462
R1388 vcc.n110 vcc.n109 1.05177
R1389 vcc.n103 vcc.n102 1.01465
R1390 vcc.n104 vcc.n24 1.00136
R1391 vcc.n143 vcc.n142 0.985286
R1392 vcc.n113 vcc.n23 0.96321
R1393 vcc.n115 vcc.n114 0.952047
R1394 vcc.n105 vcc.n103 0.936035
R1395 vcc.n131 vcc.n130 0.928261
R1396 vcc.n143 vcc.n117 0.875256
R1397 vcc.n129 vcc.n120 0.872492
R1398 vcc.n144 vcc.n143 0.862026
R1399 vcc.n109 vcc.n108 0.856347
R1400 vcc.n154 vcc.n153 0.680786
R1401 vcc.n82 vcc.n81 0.649348
R1402 vcc.n12 vcc.n3 0.492808
R1403 vcc.n130 vcc.n129 0.445398
R1404 vcc.n86 vcc.n28 0.385704
R1405 vcc.n107 vcc.n24 0.319213
R1406 vcc.n87 vcc.n86 0.283677
R1407 vcc.n153 vcc 0.255733
R1408 vcc.n82 vcc.n27 0.239152
R1409 vcc.n63 vcc.n62 0.212205
R1410 vcc.n100 vcc.n27 0.162905
R1411 vcc.n141 vcc.n140 0.137839
R1412 vcc.n130 vcc.n119 0.129667
R1413 vcc.n23 vcc.n22 0.129667
R1414 vcc.n13 vcc.n12 0.123496
R1415 vcc.n38 vcc.n25 0.114495
R1416 vcc.n85 vcc.n84 0.111978
R1417 vcc.n110 vcc.n18 0.106182
R1418 vcc.n131 vcc.n125 0.103833
R1419 vcc.n151 vcc.n150 0.0994362
R1420 vcc vcc.n154 0.0953661
R1421 vcc.n114 vcc.n109 0.09183
R1422 vcc.n152 vcc.n16 0.0866111
R1423 vcc.n56 vcc.n55 0.0819249
R1424 vcc.n105 vcc.n104 0.0791164
R1425 vcc.n86 vcc.n85 0.0730806
R1426 vcc.n106 vcc.n25 0.0728582
R1427 vcc.n87 vcc.n82 0.069878
R1428 vcc.n69 vcc.n68 0.0666499
R1429 vcc.n102 vcc 0.0571038
R1430 vcc.n70 vcc.n31 0.0501124
R1431 vcc.n132 vcc.n128 0.047375
R1432 vcc.n151 vcc.n15 0.0429528
R1433 vcc.n153 vcc.n152 0.038
R1434 vcc.n99 vcc.n28 0.0370646
R1435 vcc.n140 vcc.n118 0.0341957
R1436 vcc.n101 vcc.n100 0.0303556
R1437 vcc.n106 vcc.n105 0.0293462
R1438 vcc.n132 vcc.n131 0.0216694
R1439 vcc.n129 vcc.n118 0.020648
R1440 vcc.n54 vcc.n53 0.016785
R1441 vcc.n61 vcc.n38 0.016785
R1442 vcc.n14 vcc.n13 0.0133125
R1443 vcc.n142 vcc.n118 0.00255592
R1444 vcc.n115 vcc.n23 0.00155305
R1445 vcc.n85 vcc.n27 0.000829815
R1446 a_521_2177.n2 a_521_2177.t1 60.3532
R1447 a_521_2177.n9 a_521_2177.t3 60.3532
R1448 a_521_2177.n14 a_521_2177.n13 48.5755
R1449 a_521_2177.n0 a_521_2177.t8 19.1315
R1450 a_521_2177.n0 a_521_2177.t10 18.308
R1451 a_521_2177.n16 a_521_2177.n0 16.2724
R1452 a_521_2177.n11 a_521_2177.n10 14.6534
R1453 a_521_2177.n13 a_521_2177.t5 11.6005
R1454 a_521_2177.n13 a_521_2177.t7 11.6005
R1455 a_521_2177.n9 a_521_2177.n1 11.2227
R1456 a_521_2177.n15 a_521_2177.n14 8.08817
R1457 a_521_2177.n2 a_521_2177.n1 7.9105
R1458 a_521_2177.n3 a_521_2177.t0 3.58326
R1459 a_521_2177.n5 a_521_2177.t12 3.58326
R1460 a_521_2177.n7 a_521_2177.t15 3.58326
R1461 a_521_2177.n8 a_521_2177.t2 3.58326
R1462 a_521_2177.n3 a_521_2177.t14 3.58267
R1463 a_521_2177.n5 a_521_2177.t4 3.58267
R1464 a_521_2177.n7 a_521_2177.t6 3.58267
R1465 a_521_2177.n8 a_521_2177.t13 3.58267
R1466 a_521_2177.n12 a_521_2177.n11 3.54985
R1467 a_521_2177.n0 a_521_2177.n15 2.67636
R1468 a_521_2177.n15 a_521_2177.n1 2.10354
R1469 a_521_2177.n16 a_521_2177.t9 1.90483
R1470 a_521_2177.t11 a_521_2177.n16 1.90483
R1471 a_521_2177.n6 a_521_2177.n4 1.69798
R1472 a_521_2177.n10 a_521_2177.n8 1.61224
R1473 a_521_2177.n11 a_521_2177.n7 1.61224
R1474 a_521_2177.n6 a_521_2177.n5 1.61224
R1475 a_521_2177.n4 a_521_2177.n3 1.61224
R1476 a_521_2177.n10 a_521_2177.n9 0.995611
R1477 a_521_2177.n4 a_521_2177.n2 0.96988
R1478 a_521_2177.n14 a_521_2177.n12 0.793374
R1479 a_521_2177.n12 a_521_2177.n6 0.432312
R1480 a_8294_3178.t0 a_8294_3178.t1 53.247
R1481 vin_n.n0 vin_n.t0 21.0692
R1482 vin_n.n0 vin_n.t1 8.85313
R1483 vin_n vin_n.n0 2.40005
C0 OTA_vref_0.vb a_n832_n2063# 1.65112f
C1 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter vcc 0.512021f
C2 vin_n vin_p 2.36446f
C3 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 16.2573f
C4 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_n832_n2063# 0.002329f
C5 vcc a_1748_n2063# 0.318981f
C6 vo vcc 3.99881f
C7 vcc vin_n 0.018448f
C8 OTA_vref_0.OTA_vref_stage2_0.vref0 a_1748_n2063# 0.010991f
C9 a_458_n2063# vcc 0.335707f
C10 OTA_vref_0.OTA_vref_stage2_0.vref0 a_458_n2063# 0.011315f
C11 a_458_n2063# a_n832_n2063# 0.154422f
C12 OTA_vref_0.vb vin_n 0.374995f
C13 vcc a_3038_n2063# 0.325526f
C14 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_1748_n2063# 0.009524f
C15 OTA_vref_0.vb a_458_n2063# 3.04e-19
C16 OTA_vref_0.OTA_vref_stage2_0.vref0 a_3038_n2063# 0.112341f
C17 a_400_n1975# vcc 0.034455f
C18 OTA_vref_0.OTA_vref_stage2_0.vref0 a_400_n1975# 0.00151f
C19 a_400_n1975# a_n832_n2063# 0.10061f
C20 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_458_n2063# 0.007176f
C21 a_2980_n1975# vcc 0.034292f
C22 a_2980_n1975# OTA_vref_0.OTA_vref_stage2_0.vref0 0.037994f
C23 a_458_n2063# a_1748_n2063# 0.154516f
C24 a_400_n1975# OTA_vref_0.vb 0.036384f
C25 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_3038_n2063# 0.032619f
C26 OTA_vref_0.OTA_vref_stage2_0.vr vcc 11.4545f
C27 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter a_400_n1975# 6.62e-20
C28 a_1748_n2063# a_3038_n2063# 0.154705f
C29 OTA_vref_0.OTA_vref_stage2_0.vref0 OTA_vref_0.OTA_vref_stage2_0.vr 2.20674f
C30 OTA_vref_0.OTA_vref_stage2_0.vr a_n832_n2063# 0.369353f
C31 a_2980_n1975# OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter 0.003419f
C32 a_400_n1975# a_1748_n2063# 1.04e-19
C33 a_2980_n1975# a_1748_n2063# 0.097592f
C34 OTA_vref_0.vb OTA_vref_0.OTA_vref_stage2_0.vr 0.162898f
C35 a_400_n1975# a_458_n2063# 1.53005f
C36 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter OTA_vref_0.OTA_vref_stage2_0.vr 9.256969f
C37 OTA_vref_0.OTA_vref_stage2_0.vr a_1748_n2063# 0.341384f
C38 a_n8089_3635# vin_p 1.68092f
C39 a_2980_n1975# a_3038_n2063# 1.53765f
C40 OTA_vref_0.OTA_vref_stage2_0.vr a_458_n2063# 0.335041f
C41 a_n8089_3635# vcc 5.64e-19
C42 OTA_vref_0.OTA_vref_stage2_0.vr a_3038_n2063# 0.336282f
C43 a_400_n1975# OTA_vref_0.OTA_vref_stage2_0.vr 0.008005f
C44 OTA_vref_0.vb a_n8089_3635# 0.440922f
C45 a_2980_n1975# OTA_vref_0.OTA_vref_stage2_0.vr 0.008017f
C46 a_n8089_3635# vin_n 1.47482f
C47 vcc vin_p 0.038653f
C48 OTA_vref_0.OTA_vref_stage2_0.vref0 vcc 0.030224f
C49 vcc a_n832_n2063# 0.384127f
C50 OTA_vref_0.vb vin_p 0.158462f
C51 OTA_vref_0.vb vcc 0.288999f
C52 vo vss 10.226634f
C53 vin_n vss 14.998344f
C54 vin_p vss 14.789022f
C55 vcc vss 0.161045p
C56 OTA_vref_0.OTA_vref_stage2_0.vref0 vss 9.083215f
C57 a_2980_n1975# vss 0.471548f
C58 a_400_n1975# vss 0.471213f
C59 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter vss 25.20166f
C60 a_3038_n2063# vss 3.83372f
C61 a_1748_n2063# vss 3.70817f
C62 a_458_n2063# vss 3.70757f
C63 a_n832_n2063# vss 3.76558f
C64 OTA_vref_0.OTA_vref_stage2_0.vr vss 11.888545f
C65 OTA_vref_0.vb vss 10.2973f
C66 a_n8089_3635# vss 3.49077f
C67 vin_n.t0 vss 0.873562f
C68 vin_n.t1 vss 0.459604f
C69 vin_n.n0 vss 1.01219f
C70 a_8294_3178.t1 vss 35.8635f
C71 a_8294_3178.t0 vss 0.036479f
C72 a_521_2177.n0 vss 1.86767f
C73 a_521_2177.t9 vss 0.044291f
C74 a_521_2177.n1 vss 1.03764f
C75 a_521_2177.t1 vss 0.015632f
C76 a_521_2177.n2 vss 0.073264f
C77 a_521_2177.t0 vss 0.615961f
C78 a_521_2177.t14 vss 0.615959f
C79 a_521_2177.n3 vss 0.229584f
C80 a_521_2177.n4 vss 1.62591f
C81 a_521_2177.t12 vss 0.615961f
C82 a_521_2177.t4 vss 0.615959f
C83 a_521_2177.n5 vss 0.229584f
C84 a_521_2177.n6 vss 1.60355f
C85 a_521_2177.t15 vss 0.615961f
C86 a_521_2177.t6 vss 0.615959f
C87 a_521_2177.n7 vss 0.229584f
C88 a_521_2177.t2 vss 0.615961f
C89 a_521_2177.t13 vss 0.615959f
C90 a_521_2177.n8 vss 0.229584f
C91 a_521_2177.t3 vss 0.015632f
C92 a_521_2177.n9 vss 0.202745f
C93 a_521_2177.n10 vss 1.62929f
C94 a_521_2177.n11 vss 1.6494f
C95 a_521_2177.n12 vss 0.10423f
C96 a_521_2177.t5 vss 0.004429f
C97 a_521_2177.t7 vss 0.004429f
C98 a_521_2177.n13 vss 0.009369f
C99 a_521_2177.n14 vss 0.034107f
C100 a_521_2177.n15 vss 0.623005f
C101 a_521_2177.t10 vss 0.202079f
C102 a_521_2177.t8 vss 0.223388f
C103 a_521_2177.n16 vss 0.139622f
C104 a_521_2177.t11 vss 0.044291f
C105 vcc.t23 vss 0.004163f
C106 vcc.t26 vss 0.004163f
C107 vcc.n0 vss 0.009136f
C108 vcc.t24 vss 0.004163f
C109 vcc.t27 vss 0.004163f
C110 vcc.n1 vss 0.008699f
C111 vcc.n2 vss 0.09654f
C112 vcc.n3 vss 0.645547f
C113 vcc.n4 vss 0.46291f
C114 vcc.n5 vss 0.123276f
C115 vcc.n6 vss 0.123276f
C116 vcc.n7 vss 0.849849f
C117 vcc.n8 vss 1.46396f
C118 vcc.t22 vss 2.29696f
C119 vcc.n9 vss 2.15172f
C120 vcc.t25 vss 2.29666f
C121 vcc.n10 vss 1.46191f
C122 vcc.n11 vss 0.915581f
C123 vcc.n12 vss 0.81811f
C124 vcc.n13 vss 1.09885f
C125 vcc.n14 vss 0.74524f
C126 vcc.n15 vss 0.676498f
C127 vcc.n16 vss 0.427825f
C128 vcc.n17 vss 0.283327f
C129 vcc.n18 vss 0.347517f
C130 vcc.n19 vss 0.13567f
C131 vcc.n20 vss 0.135643f
C132 vcc.n21 vss 0.618633f
C133 vcc.n22 vss 0.00533f
C134 vcc.n23 vss 0.079017f
C135 vcc.t15 vss 0.00867f
C136 vcc.t11 vss 0.008671f
C137 vcc.n24 vss 0.141204f
C138 vcc.n25 vss 0.093082f
C139 vcc.t3 vss 0.008671f
C140 vcc.t9 vss 0.008671f
C141 vcc.t5 vss 0.002313f
C142 vcc.t13 vss 0.002313f
C143 vcc.n26 vss 0.004934f
C144 vcc.n27 vss 0.25323f
C145 vcc.n28 vss 0.029076f
C146 vcc.n29 vss 0.081294f
C147 vcc.n30 vss 0.025909f
C148 vcc.n31 vss 0.071257f
C149 vcc.n32 vss 0.124324f
C150 vcc.n33 vss 0.124324f
C151 vcc.n34 vss 0.028041f
C152 vcc.n35 vss 0.111776f
C153 vcc.n37 vss 0.016442f
C154 vcc.n38 vss 0.019888f
C155 vcc.n40 vss 0.029982f
C156 vcc.n41 vss 0.016442f
C157 vcc.n42 vss 0.109561f
C158 vcc.n43 vss 0.030548f
C159 vcc.n44 vss 0.360105f
C160 vcc.n45 vss 0.023657f
C161 vcc.n46 vss 0.023657f
C162 vcc.n47 vss 0.047455f
C163 vcc.n48 vss 0.101104f
C164 vcc.n49 vss 0.135092f
C165 vcc.t14 vss 0.16502f
C166 vcc.n50 vss 0.147129f
C167 vcc.t10 vss 0.16497f
C168 vcc.n51 vss 0.131328f
C169 vcc.n52 vss 0.015722f
C170 vcc.n53 vss 0.061827f
C171 vcc.n54 vss 0.174973f
C172 vcc.n55 vss 0.19442f
C173 vcc.n56 vss 0.074644f
C174 vcc.n57 vss 0.124324f
C175 vcc.t16 vss 0.187548f
C176 vcc.n59 vss 0.016442f
C177 vcc.n60 vss 0.124324f
C178 vcc.n61 vss 0.185565f
C179 vcc.n62 vss 0.205026f
C180 vcc.n63 vss 0.071707f
C181 vcc.n64 vss 0.124324f
C182 vcc.t2 vss 0.187548f
C183 vcc.n66 vss 0.016442f
C184 vcc.n67 vss 0.124324f
C185 vcc.n68 vss 0.072221f
C186 vcc.n69 vss 0.201829f
C187 vcc.n70 vss 0.200423f
C188 vcc.n71 vss 0.029301f
C189 vcc.n72 vss 0.016442f
C190 vcc.t8 vss 0.187548f
C191 vcc.n75 vss 0.016442f
C192 vcc.n76 vss 0.113787f
C193 vcc.n77 vss 0.13533f
C194 vcc.n78 vss 0.027286f
C195 vcc.n79 vss 0.048891f
C196 vcc.t12 vss 0.092818f
C197 vcc.n80 vss 0.154676f
C198 vcc.n81 vss 0.078226f
C199 vcc.n82 vss 0.086197f
C200 vcc.t1 vss 0.001157f
C201 vcc.t7 vss 0.001157f
C202 vcc.n83 vss 0.002423f
C203 vcc.n84 vss 0.26556f
C204 vcc.n85 vss 0.051237f
C205 vcc.n86 vss 0.14154f
C206 vcc.n87 vss 0.338875f
C207 vcc.n88 vss 0.04544f
C208 vcc.n89 vss 0.03647f
C209 vcc.t0 vss 0.192908f
C210 vcc.t4 vss 0.174646f
C211 vcc.n90 vss 0.143103f
C212 vcc.t6 vss 0.061595f
C213 vcc.n91 vss 0.115617f
C214 vcc.n92 vss 0.03647f
C215 vcc.n93 vss 0.027286f
C216 vcc.n94 vss 0.042735f
C217 vcc.n95 vss 0.112946f
C218 vcc.n96 vss 0.013544f
C219 vcc.n97 vss 0.153098f
C220 vcc.n98 vss 0.086093f
C221 vcc.n99 vss 0.06173f
C222 vcc.n100 vss 0.089038f
C223 vcc.n101 vss 0.159668f
C224 vcc.n102 vss 0.113163f
C225 vcc.n103 vss 0.184054f
C226 vcc.t17 vss 0.008671f
C227 vcc.n104 vss 0.114258f
C228 vcc.n105 vss 0.081797f
C229 vcc.n106 vss 0.507191f
C230 vcc.n107 vss 0.113621f
C231 vcc.n108 vss 1.17528f
C232 vcc.n109 vss 1.52141f
C233 vcc.n110 vss 0.571893f
C234 vcc.n111 vss 0.077213f
C235 vcc.n112 vss 0.246651f
C236 vcc.n113 vss 0.193519f
C237 vcc.n114 vss 0.151016f
C238 vcc.n115 vss 0.388432f
C239 vcc.n116 vss 0.146777f
C240 vcc.n117 vss 0.488438f
C241 vcc.n118 vss 0.006547f
C242 vcc.n119 vss 0.112248f
C243 vcc.n120 vss 1.56005f
C244 vcc.n121 vss 0.34927f
C245 vcc.n122 vss 0.34927f
C246 vcc.t30 vss 0.557597f
C247 vcc.t28 vss 0.459583f
C248 vcc.n123 vss 0.380591f
C249 vcc.n124 vss 0.262255f
C250 vcc.n125 vss 0.216741f
C251 vcc.t31 vss 0.016191f
C252 vcc.t29 vss 0.016191f
C253 vcc.n126 vss 0.042058f
C254 vcc.t35 vss 0.016191f
C255 vcc.t33 vss 0.016191f
C256 vcc.n127 vss 0.041282f
C257 vcc.n128 vss 0.660578f
C258 vcc.n129 vss 1.12219f
C259 vcc.n130 vss 0.276206f
C260 vcc.n131 vss 0.19639f
C261 vcc.n132 vss 0.21066f
C262 vcc.n133 vss 0.01607f
C263 vcc.n134 vss 0.237598f
C264 vcc.n135 vss 0.049221f
C265 vcc.t32 vss 0.557597f
C266 vcc.t34 vss 0.459583f
C267 vcc.n136 vss 0.306389f
C268 vcc.n137 vss 0.049221f
C269 vcc.n138 vss 0.572378f
C270 vcc.n139 vss 0.322156f
C271 vcc.n140 vss 0.011894f
C272 vcc.n141 vss 0.444899f
C273 vcc.n142 vss 0.290962f
C274 vcc.n143 vss 0.44643f
C275 vcc.n144 vss 0.203314f
C276 vcc.n145 vss 0.614715f
C277 vcc.n146 vss 2.68269f
C278 vcc.t18 vss 3.17686f
C279 vcc.t21 vss 1.89988f
C280 vcc.n147 vss 1.35529f
C281 vcc.t19 vss 2.16598f
C282 vcc.t20 vss 2.90944f
C283 vcc.n148 vss 2.25081f
C284 vcc.n149 vss 0.383538f
C285 vcc.n150 vss 0.463313f
C286 vcc.n151 vss 0.468512f
C287 vcc.n152 vss 0.480372f
C288 vcc.n153 vss 0.930633f
C289 vcc.n154 vss 0.22892f
C290 a_959_2177.t4 vss 0.216942f
C291 a_959_2177.t0 vss 0.216942f
C292 a_959_2177.t5 vss 0.216942f
C293 a_959_2177.n0 vss 0.671366f
C294 a_959_2177.t6 vss 0.216942f
C295 a_959_2177.t2 vss 0.216942f
C296 a_959_2177.n1 vss 0.762068f
C297 a_959_2177.n2 vss 4.7253f
C298 a_959_2177.t8 vss 0.399519f
C299 a_959_2177.t9 vss 0.10124f
C300 a_959_2177.t10 vss 0.10124f
C301 a_959_2177.n3 vss 0.235864f
C302 a_959_2177.t11 vss 0.427351f
C303 a_959_2177.n4 vss 2.07187f
C304 a_959_2177.n5 vss 1.4064f
C305 a_959_2177.n6 vss 2.8881f
C306 a_959_2177.t1 vss 0.216942f
C307 a_959_2177.t7 vss 0.216942f
C308 a_959_2177.n7 vss 0.76209f
C309 a_959_2177.n8 vss 3.54056f
C310 a_959_2177.n9 vss 0.671495f
C311 a_959_2177.t3 vss 0.216942f
C312 vo.t5 vss 0.100527f
C313 vo.t2 vss 0.737707f
C314 vo.t3 vss 0.8199f
C315 vo.n0 vss 4.30681f
C316 vo.t1 vss 0.155102f
C317 vo.t4 vss 0.155102f
C318 vo.n1 vss 0.430799f
C319 vo.n2 vss 2.50099f
C320 vo.t7 vss 0.084327f
C321 vo.n3 vss 2.47737f
C322 vo.t8 vss 0.076075f
C323 vo.n4 vss 1.14312f
C324 vo.n5 vss 0.767691f
C325 vo.t6 vss 0.01551f
C326 vo.t0 vss 0.01551f
C327 vo.n6 vss 0.090416f
C328 vo.n7 vss 2.00431f
C329 OTA_stage2_0.vd1.n0 vss 18.8388f
C330 OTA_stage2_0.vd1.t2 vss 37.7439f
C331 OTA_stage2_0.vd1.t8 vss 1.71875f
C332 OTA_stage2_0.vd1.t5 vss 1.73013f
C333 OTA_stage2_0.vd1.t7 vss 1.73013f
C334 OTA_stage2_0.vd1.t6 vss 1.71875f
C335 OTA_stage2_0.vd1.t4 vss 0.046875f
C336 OTA_stage2_0.vd1.t3 vss 0.051839f
C337 OTA_stage2_0.vd1.t0 vss 0.385333f
C338 OTA_stage2_0.vd1.t1 vss 0.235537f
C339 OTA_vref_0.vb1.n0 vss 5.67164f
C340 OTA_vref_0.vb1.n1 vss 0.347123f
C341 OTA_vref_0.OTA_vref_stage2_0.vb1 vss 1.42021f
C342 OTA_vref_0.vb1.t7 vss 0.8461f
C343 OTA_vref_0.vb1.t6 vss 0.834437f
C344 OTA_vref_0.vb1.t9 vss 0.834437f
C345 OTA_vref_0.vb1.t8 vss 0.834437f
C346 OTA_stage2_0.vb1 vss 0.916273f
C347 OTA_vref_0.vb1.t2 vss 0.006934f
C348 OTA_vref_0.vb1.t5 vss 0.006934f
C349 OTA_vref_0.vb1.n2 vss 0.018589f
C350 OTA_vref_0.vb1.t1 vss 0.006934f
C351 OTA_vref_0.vb1.t0 vss 0.006934f
C352 OTA_vref_0.vb1.n3 vss 0.017571f
C353 OTA_vref_0.vb1.t4 vss 0.006934f
C354 OTA_vref_0.vb1.t3 vss 0.006934f
C355 OTA_vref_0.vb1.n4 vss 0.017571f
C356 OTA_stage2_0.vd2.t0 vss 39.2136f
C357 OTA_stage2_0.vd2.t4 vss 1.3368f
C358 OTA_stage2_0.vd2.t5 vss 1.33009f
C359 OTA_stage2_0.vd2.t3 vss 1.33009f
C360 OTA_stage2_0.vd2.t6 vss 1.32145f
C361 OTA_stage2_0.vd2.t2 vss 0.033976f
C362 OTA_stage2_0.vd2.t1 vss 0.033964f
C363 vin_p.t0 vss 0.87648f
C364 vin_p.t1 vss 0.460642f
C365 vin_p.n0 vss 1.00726f
C366 OTA_vref_0.OTA_vref_stage2_0.vr.t22 vss 0.304639f
C367 OTA_vref_0.OTA_vref_stage2_0.vr.t25 vss 0.304639f
C368 OTA_vref_0.OTA_vref_stage2_0.vr.t1 vss 0.025938f
C369 OTA_vref_0.OTA_vref_stage2_0.vr.t3 vss 0.025974f
C370 OTA_vref_0.OTA_vref_stage2_0.vr.t2 vss 0.460559f
C371 OTA_vref_0.OTA_vref_stage2_0.vr.n0 vss 0.83568f
C372 OTA_vref_0.OTA_vref_stage2_0.vr.t10 vss 0.277156f
C373 OTA_vref_0.OTA_vref_stage2_0.vr.t9 vss 0.054965f
C374 OTA_vref_0.OTA_vref_stage2_0.vr.t14 vss 0.054965f
C375 OTA_vref_0.OTA_vref_stage2_0.vr.n1 vss 0.208795f
C376 OTA_vref_0.OTA_vref_stage2_0.vr.t11 vss 0.054965f
C377 OTA_vref_0.OTA_vref_stage2_0.vr.t16 vss 0.054965f
C378 OTA_vref_0.OTA_vref_stage2_0.vr.n2 vss 0.208795f
C379 OTA_vref_0.OTA_vref_stage2_0.vr.t13 vss 0.054965f
C380 OTA_vref_0.OTA_vref_stage2_0.vr.t6 vss 0.054965f
C381 OTA_vref_0.OTA_vref_stage2_0.vr.n3 vss 0.208795f
C382 OTA_vref_0.OTA_vref_stage2_0.vr.t8 vss 0.302577f
C383 OTA_vref_0.OTA_vref_stage2_0.vr.n4 vss 1.71656f
C384 OTA_vref_0.OTA_vref_stage2_0.vr.n5 vss 0.983628f
C385 OTA_vref_0.OTA_vref_stage2_0.vr.n6 vss 0.983628f
C386 OTA_vref_0.OTA_vref_stage2_0.vr.n7 vss 0.924068f
C387 OTA_vref_0.OTA_vref_stage2_0.vr.t15 vss 0.054965f
C388 OTA_vref_0.OTA_vref_stage2_0.vr.t7 vss 0.054965f
C389 OTA_vref_0.OTA_vref_stage2_0.vr.n8 vss 0.208795f
C390 OTA_vref_0.OTA_vref_stage2_0.vr.t4 vss 0.054965f
C391 OTA_vref_0.OTA_vref_stage2_0.vr.t18 vss 0.054965f
C392 OTA_vref_0.OTA_vref_stage2_0.vr.n9 vss 0.208795f
C393 OTA_vref_0.OTA_vref_stage2_0.vr.t12 vss 0.054965f
C394 OTA_vref_0.OTA_vref_stage2_0.vr.t5 vss 0.054965f
C395 OTA_vref_0.OTA_vref_stage2_0.vr.n10 vss 0.23714f
C396 OTA_vref_0.OTA_vref_stage2_0.vr.n11 vss 1.67206f
C397 OTA_vref_0.OTA_vref_stage2_0.vr.n12 vss 0.983628f
C398 OTA_vref_0.OTA_vref_stage2_0.vr.t19 vss 0.054965f
C399 OTA_vref_0.OTA_vref_stage2_0.vr.t17 vss 0.054965f
C400 OTA_vref_0.OTA_vref_stage2_0.vr.n13 vss 0.208795f
C401 OTA_vref_0.OTA_vref_stage2_0.vr.n14 vss 1.02084f
C402 OTA_vref_0.OTA_vref_stage2_0.vr.n15 vss 1.69107f
C403 OTA_vref_0.OTA_vref_stage2_0.vr.n16 vss 0.847025f
C404 OTA_vref_0.OTA_vref_stage2_0.vr.t0 vss 0.460559f
C405 OTA_vref_0.OTA_vref_stage2_0.vr.n17 vss 0.780032f
C406 OTA_vref_0.OTA_vref_stage2_0.vr.n18 vss 0.111572f
C407 OTA_vref_0.OTA_vref_stage2_0.vr.n19 vss 0.371836f
C408 OTA_vref_0.OTA_vref_stage2_0.vr.n20 vss 0.367258f
C409 OTA_vref_0.OTA_vref_stage2_0.vr.t21 vss 0.610236f
C410 OTA_vref_0.OTA_vref_stage2_0.vr.t23 vss 0.586815f
C411 OTA_vref_0.OTA_vref_stage2_0.vr.n21 vss 1.65918f
C412 OTA_vref_0.OTA_vref_stage2_0.vr.t20 vss 0.586815f
C413 OTA_vref_0.OTA_vref_stage2_0.vr.n22 vss 0.980201f
C414 OTA_vref_0.OTA_vref_stage2_0.vr.t26 vss 0.586815f
C415 OTA_vref_0.OTA_vref_stage2_0.vr.n23 vss 0.978893f
C416 OTA_vref_0.OTA_vref_stage2_0.vr.t24 vss 0.586815f
C417 OTA_vref_0.OTA_vref_stage2_0.vr.n24 vss 0.894432f
C418 OTA_vref_0.OTA_vref_stage2_0.vref0.n0 vss 1.12775f
C419 OTA_vref_0.OTA_vref_stage2_0.vref0.t32 vss 0.077096f
C420 OTA_vref_0.OTA_vref_stage2_0.vref0.t3 vss 0.07938f
C421 OTA_vref_0.OTA_vref_stage2_0.vref0.t7 vss 0.07938f
C422 OTA_vref_0.OTA_vref_stage2_0.vref0.n1 vss 0.254851f
C423 OTA_vref_0.OTA_vref_stage2_0.vref0.t11 vss 0.07938f
C424 OTA_vref_0.OTA_vref_stage2_0.vref0.t24 vss 0.07938f
C425 OTA_vref_0.OTA_vref_stage2_0.vref0.n2 vss 0.254735f
C426 OTA_vref_0.OTA_vref_stage2_0.vref0.t16 vss 0.07938f
C427 OTA_vref_0.OTA_vref_stage2_0.vref0.t1 vss 0.07938f
C428 OTA_vref_0.OTA_vref_stage2_0.vref0.n3 vss 0.278086f
C429 OTA_vref_0.OTA_vref_stage2_0.vref0.t29 vss 0.07938f
C430 OTA_vref_0.OTA_vref_stage2_0.vref0.t20 vss 0.07938f
C431 OTA_vref_0.OTA_vref_stage2_0.vref0.n4 vss 0.254416f
C432 OTA_vref_0.OTA_vref_stage2_0.vref0.n5 vss 1.7151f
C433 OTA_vref_0.OTA_vref_stage2_0.vref0.t13 vss 0.07938f
C434 OTA_vref_0.OTA_vref_stage2_0.vref0.t0 vss 0.07938f
C435 OTA_vref_0.OTA_vref_stage2_0.vref0.n6 vss 0.254416f
C436 OTA_vref_0.OTA_vref_stage2_0.vref0.n7 vss 0.92465f
C437 OTA_vref_0.OTA_vref_stage2_0.vref0.t26 vss 0.07938f
C438 OTA_vref_0.OTA_vref_stage2_0.vref0.t6 vss 0.07938f
C439 OTA_vref_0.OTA_vref_stage2_0.vref0.n8 vss 0.254416f
C440 OTA_vref_0.OTA_vref_stage2_0.vref0.n9 vss 0.92465f
C441 OTA_vref_0.OTA_vref_stage2_0.vref0.t10 vss 0.07938f
C442 OTA_vref_0.OTA_vref_stage2_0.vref0.t21 vss 0.07938f
C443 OTA_vref_0.OTA_vref_stage2_0.vref0.n10 vss 0.254416f
C444 OTA_vref_0.OTA_vref_stage2_0.vref0.n11 vss 0.92465f
C445 OTA_vref_0.OTA_vref_stage2_0.vref0.t4 vss 0.07938f
C446 OTA_vref_0.OTA_vref_stage2_0.vref0.t19 vss 0.07938f
C447 OTA_vref_0.OTA_vref_stage2_0.vref0.n12 vss 0.254416f
C448 OTA_vref_0.OTA_vref_stage2_0.vref0.n13 vss 0.92465f
C449 OTA_vref_0.OTA_vref_stage2_0.vref0.t12 vss 0.07938f
C450 OTA_vref_0.OTA_vref_stage2_0.vref0.t23 vss 0.07938f
C451 OTA_vref_0.OTA_vref_stage2_0.vref0.n14 vss 0.254416f
C452 OTA_vref_0.OTA_vref_stage2_0.vref0.n15 vss 0.92465f
C453 OTA_vref_0.OTA_vref_stage2_0.vref0.t22 vss 0.07938f
C454 OTA_vref_0.OTA_vref_stage2_0.vref0.t18 vss 0.07938f
C455 OTA_vref_0.OTA_vref_stage2_0.vref0.n16 vss 0.254416f
C456 OTA_vref_0.OTA_vref_stage2_0.vref0.n17 vss 1.43858f
C457 OTA_vref_0.OTA_vref_stage2_0.vref0.n18 vss 1.30683f
C458 OTA_vref_0.OTA_vref_stage2_0.vref0.t14 vss 0.07938f
C459 OTA_vref_0.OTA_vref_stage2_0.vref0.t27 vss 0.07938f
C460 OTA_vref_0.OTA_vref_stage2_0.vref0.n19 vss 0.254851f
C461 OTA_vref_0.OTA_vref_stage2_0.vref0.t2 vss 0.07938f
C462 OTA_vref_0.OTA_vref_stage2_0.vref0.t5 vss 0.07938f
C463 OTA_vref_0.OTA_vref_stage2_0.vref0.n20 vss 0.254851f
C464 OTA_vref_0.OTA_vref_stage2_0.vref0.t17 vss 0.07938f
C465 OTA_vref_0.OTA_vref_stage2_0.vref0.t31 vss 0.07938f
C466 OTA_vref_0.OTA_vref_stage2_0.vref0.n21 vss 0.254851f
C467 OTA_vref_0.OTA_vref_stage2_0.vref0.t25 vss 0.07938f
C468 OTA_vref_0.OTA_vref_stage2_0.vref0.t8 vss 0.07938f
C469 OTA_vref_0.OTA_vref_stage2_0.vref0.n22 vss 0.254851f
C470 OTA_vref_0.OTA_vref_stage2_0.vref0.t15 vss 0.07938f
C471 OTA_vref_0.OTA_vref_stage2_0.vref0.t28 vss 0.07938f
C472 OTA_vref_0.OTA_vref_stage2_0.vref0.n23 vss 0.254851f
C473 OTA_vref_0.OTA_vref_stage2_0.vref0.t30 vss 0.07938f
C474 OTA_vref_0.OTA_vref_stage2_0.vref0.t9 vss 0.07938f
C475 OTA_vref_0.OTA_vref_stage2_0.vref0.n24 vss 0.264844f
C476 OTA_vref_0.OTA_vref_stage2_0.vref0.n25 vss 1.60894f
C477 OTA_vref_0.OTA_vref_stage2_0.vref0.n26 vss 0.933767f
C478 OTA_vref_0.OTA_vref_stage2_0.vref0.n27 vss 0.933767f
C479 OTA_vref_0.OTA_vref_stage2_0.vref0.n28 vss 0.933767f
C480 OTA_vref_0.OTA_vref_stage2_0.vref0.n29 vss 0.914004f
C481 a_n27_n4200.n0 vss 0.646091f
C482 a_n27_n4200.n1 vss 0.42162f
C483 a_n27_n4200.n2 vss 0.651883f
C484 a_n27_n4200.n3 vss 0.42562f
C485 a_n27_n4200.n4 vss 0.434861f
C486 a_n27_n4200.n6 vss 0.527809f
C487 a_n27_n4200.n7 vss 0.058555f
C488 a_n27_n4200.n9 vss 0.564683f
C489 a_n27_n4200.n10 vss 0.06018f
C490 a_n27_n4200.n11 vss 0.06069f
C491 a_n27_n4200.n12 vss 0.564177f
C492 a_n27_n4200.n14 vss 0.450822f
C493 a_n27_n4200.n16 vss 0.543856f
C494 a_n27_n4200.n17 vss 0.063412f
C495 a_n27_n4200.n18 vss 0.569986f
C496 a_n27_n4200.n20 vss 0.589474f
C497 a_n27_n4200.n21 vss 0.875998f
C498 a_n27_n4200.n22 vss 0.414104f
C499 a_n27_n4200.n23 vss 0.598858f
C500 a_n27_n4200.n24 vss 0.589368f
C501 a_n27_n4200.n25 vss 0.751854f
C502 a_n27_n4200.n26 vss 0.589533f
C503 a_n27_n4200.n27 vss 0.589369f
C504 a_n27_n4200.n28 vss 0.279618f
C505 a_n27_n4200.n30 vss 0.592443f
C506 a_n27_n4200.n31 vss 0.283642f
C507 a_n27_n4200.n32 vss 0.233813f
C508 a_n27_n4200.n33 vss 0.447151f
C509 a_n27_n4200.n34 vss 0.447748f
C510 a_n27_n4200.t30 vss 0.426145f
C511 a_n27_n4200.t26 vss 0.426145f
C512 a_n27_n4200.n35 vss 0.159721f
C513 a_n27_n4200.t34 vss 0.036484f
C514 a_n27_n4200.t25 vss 0.036484f
C515 a_n27_n4200.t43 vss 0.036484f
C516 a_n27_n4200.n36 vss 0.077937f
C517 a_n27_n4200.t24 vss 0.426781f
C518 a_n27_n4200.n37 vss 0.509606f
C519 a_n27_n4200.t46 vss 0.036484f
C520 a_n27_n4200.t15 vss 0.036484f
C521 a_n27_n4200.n38 vss 0.078094f
C522 a_n27_n4200.t14 vss 0.427925f
C523 a_n27_n4200.t22 vss 0.426145f
C524 a_n27_n4200.t23 vss 0.036484f
C525 a_n27_n4200.t42 vss 0.036484f
C526 a_n27_n4200.n39 vss 0.077885f
C527 a_n27_n4200.t45 vss 0.036484f
C528 a_n27_n4200.t13 vss 0.036484f
C529 a_n27_n4200.n40 vss 0.077885f
C530 a_n27_n4200.t6 vss 0.426145f
C531 a_n27_n4200.t31 vss 0.036484f
C532 a_n27_n4200.t40 vss 0.036484f
C533 a_n27_n4200.n41 vss 0.077937f
C534 a_n27_n4200.t36 vss 0.036484f
C535 a_n27_n4200.t9 vss 0.036484f
C536 a_n27_n4200.n42 vss 0.077937f
C537 a_n27_n4200.t8 vss 0.426145f
C538 a_n27_n4200.t28 vss 0.426145f
C539 a_n27_n4200.t29 vss 0.036484f
C540 a_n27_n4200.t44 vss 0.036484f
C541 a_n27_n4200.n43 vss 0.077939f
C542 a_n27_n4200.t33 vss 0.036484f
C543 a_n27_n4200.t19 vss 0.036484f
C544 a_n27_n4200.n44 vss 0.077937f
C545 a_n27_n4200.t18 vss 0.426145f
C546 a_n27_n4200.t21 vss 0.036484f
C547 a_n27_n4200.t41 vss 0.036484f
C548 a_n27_n4200.n45 vss 0.077885f
C549 a_n27_n4200.t47 vss 0.036484f
C550 a_n27_n4200.t17 vss 0.036484f
C551 a_n27_n4200.n46 vss 0.077885f
C552 a_n27_n4200.t16 vss 0.426145f
C553 a_n27_n4200.t4 vss 0.426145f
C554 a_n27_n4200.t5 vss 0.036484f
C555 a_n27_n4200.t38 vss 0.036484f
C556 a_n27_n4200.n47 vss 0.077885f
C557 a_n27_n4200.t10 vss 0.426788f
C558 a_n27_n4200.n48 vss 0.499272f
C559 a_n27_n4200.t37 vss 0.036484f
C560 a_n27_n4200.t11 vss 0.036484f
C561 a_n27_n4200.n49 vss 0.077937f
C562 a_n27_n4200.t27 vss 0.036484f
C563 a_n27_n4200.t39 vss 0.036484f
C564 a_n27_n4200.n50 vss 0.077937f
C565 a_n27_n4200.n51 vss 0.1597f
C566 a_n27_n4200.n52 vss 0.173683f
C567 a_n27_n4200.t20 vss 0.426145f
C568 a_n27_n4200.t35 vss 0.036484f
C569 a_n27_n4200.t7 vss 0.036484f
C570 a_n27_n4200.n53 vss 0.077885f
C571 a_n27_n4200.t3 vss 0.036484f
C572 a_n27_n4200.t32 vss 0.036484f
C573 a_n27_n4200.n54 vss 0.077885f
C574 a_n27_n4200.t12 vss 0.427916f
C575 a_n27_n4200.t2 vss 0.426145f
C576 a_n27_n4200.n55 vss 0.173683f
C577 a_n27_n4200.n56 vss 0.1597f
C578 a_n27_n4200.t0 vss 0.426145f
C579 a_n27_n4200.n57 vss 0.077937f
C580 a_n27_n4200.t1 vss 0.036484f
C581 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n0 vss 0.108958f
C582 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n1 vss 0.122425f
C583 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n2 vss 0.215214f
C584 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t0 vss 0.10796f
C585 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n3 vss 0.122425f
C586 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t24 vss 0.478982f
C587 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t16 vss 0.480213f
C588 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n4 vss 1.17119f
C589 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n5 vss 0.305431f
C590 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t17 vss 0.478883f
C591 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n6 vss 0.233332f
C592 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n7 vss 0.470573f
C593 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t13 vss 0.478028f
C594 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n8 vss 0.470573f
C595 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t32 vss 0.478028f
C596 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n10 vss 0.470128f
C597 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t26 vss 0.478028f
C598 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n11 vss 0.119324f
C599 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n12 vss 0.391163f
C600 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n13 vss 0.207747f
C601 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n14 vss 0.305316f
C602 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t19 vss 0.478028f
C603 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n15 vss 0.222808f
C604 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n16 vss 0.474153f
C605 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t12 vss 0.478028f
C606 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n18 vss 0.474153f
C607 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t31 vss 0.478028f
C608 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n20 vss 0.472108f
C609 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t3 vss 0.478028f
C610 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n21 vss 0.114608f
C611 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n22 vss 0.358069f
C612 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n23 vss 0.171291f
C613 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n24 vss 0.305164f
C614 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t14 vss 0.478885f
C615 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n25 vss 0.233869f
C616 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n26 vss 0.471116f
C617 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t34 vss 0.478028f
C618 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n27 vss 0.471116f
C619 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t5 vss 0.478028f
C620 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n29 vss 0.471016f
C621 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t27 vss 0.478028f
C622 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n30 vss 0.116651f
C623 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n31 vss 0.391917f
C624 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n32 vss 0.175402f
C625 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n33 vss 0.305187f
C626 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t25 vss 0.478028f
C627 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n34 vss 0.233649f
C628 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n35 vss 0.470031f
C629 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t15 vss 0.478028f
C630 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n37 vss 0.470031f
C631 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t9 vss 0.478028f
C632 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n39 vss 0.470335f
C633 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t29 vss 0.478028f
C634 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n40 vss 0.118954f
C635 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n41 vss 0.357235f
C636 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n42 vss 0.171379f
C637 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n43 vss 0.305728f
C638 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t18 vss 0.478865f
C639 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n44 vss 0.230684f
C640 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n45 vss 0.470852f
C641 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t10 vss 0.478028f
C642 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n46 vss 0.470852f
C643 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t30 vss 0.478028f
C644 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n48 vss 0.466741f
C645 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t33 vss 0.478028f
C646 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n49 vss 0.124091f
C647 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n50 vss 0.391922f
C648 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n51 vss 0.175402f
C649 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t6 vss 0.478028f
C650 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n52 vss 0.282661f
C651 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n53 vss 0.46793f
C652 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t21 vss 0.478926f
C653 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n54 vss 0.239387f
C654 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t22 vss 0.478028f
C655 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n55 vss 0.46793f
C656 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n56 vss 0.304748f
C657 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t11 vss 0.478028f
C658 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n58 vss 0.303873f
C659 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n59 vss 0.15773f
C660 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n60 vss 0.205168f
C661 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n61 vss 0.171854f
C662 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n62 vss 0.305508f
C663 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t23 vss 0.478842f
C664 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n63 vss 0.227626f
C665 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n64 vss 0.473853f
C666 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t4 vss 0.478028f
C667 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n65 vss 0.473853f
C668 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t7 vss 0.478028f
C669 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n67 vss 0.473079f
C670 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t28 vss 0.478028f
C671 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n68 vss 0.113695f
C672 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n69 vss 0.395354f
C673 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n70 vss 0.17643f
C674 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t8 vss 0.478987f
C675 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t20 vss 0.480409f
C676 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n71 vss 1.18521f
C677 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n72 vss 0.383032f
C678 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n73 vss 0.604284f
C679 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n74 vss 0.490623f
C680 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n75 vss 0.45162f
C681 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n76 vss 0.184059f
C682 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n77 vss 0.215214f
C683 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n78 vss 0.215214f
C684 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n79 vss 0.110183f
C685 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n80 vss 0.110183f
C686 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n81 vss 0.122425f
C687 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n82 vss 0.109159f
C688 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n83 vss 0.21592f
C689 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n84 vss 0.21592f
C690 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n85 vss -6.43681f
C691 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n86 vss 6.71166f
C692 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n87 vss 0.329447f
C693 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t2 vss 0.041255f
C694 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.t1 vss 0.04125f
C695 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n88 vss 1.0567f
C696 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n89 vss 0.591984f
C697 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n90 vss 0.201225f
C698 OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter.n91 vss 0.059988f
.ends

