VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DalinEM_diff_amp
  CLASS BLOCK ;
  FOREIGN tt_um_DalinEM_diff_amp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 14.355000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.524000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 288.000000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 288.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 15.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 170.201599 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 157.000 5.000 159.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.000 5.000 4.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 43.815 130.925 83.865 138.300 ;
      LAYER pwell ;
        RECT 43.835 113.355 48.935 120.315 ;
        RECT 50.135 110.700 77.770 128.475 ;
        RECT 50.555 110.530 50.670 110.700 ;
        RECT 51.140 110.530 77.305 110.540 ;
      LAYER nwell ;
        RECT 86.210 110.535 99.275 149.330 ;
        RECT 111.390 111.180 121.420 120.370 ;
      LAYER pwell ;
        RECT 125.970 113.220 127.980 120.040 ;
      LAYER nwell ;
        RECT 79.835 94.205 86.700 97.380 ;
        RECT 107.550 97.315 117.605 97.320 ;
        RECT 89.220 94.125 93.180 97.315 ;
        RECT 95.670 94.125 99.630 97.315 ;
        RECT 102.120 94.125 106.080 97.315 ;
        RECT 107.550 94.160 117.625 97.315 ;
        RECT 111.705 94.155 117.625 94.160 ;
      LAYER pwell ;
        RECT 79.765 89.665 108.135 93.900 ;
        RECT 110.725 92.850 117.425 93.615 ;
        RECT 110.725 87.680 111.490 92.850 ;
        RECT 116.660 87.680 117.425 92.850 ;
        RECT 110.725 86.915 117.425 87.680 ;
        RECT 83.485 77.600 117.695 86.685 ;
        RECT 83.485 77.585 106.740 77.600 ;
        RECT 106.905 77.585 117.695 77.600 ;
        RECT 83.485 77.355 117.695 77.585 ;
        RECT 83.485 77.335 106.735 77.355 ;
        RECT 106.895 77.335 117.695 77.355 ;
        RECT 83.485 71.115 117.695 77.335 ;
        RECT 13.425 41.735 28.995 52.525 ;
      LAYER nwell ;
        RECT 36.465 52.435 39.625 52.455 ;
      LAYER pwell ;
        RECT 29.225 51.490 35.925 52.255 ;
        RECT 29.225 46.320 29.990 51.490 ;
        RECT 35.160 46.320 35.925 51.490 ;
      LAYER nwell ;
        RECT 36.465 46.535 39.630 52.435 ;
        RECT 89.160 47.705 129.210 55.080 ;
      LAYER pwell ;
        RECT 29.225 45.555 35.925 46.320 ;
        RECT 13.425 41.725 19.895 41.735 ;
        RECT 13.425 41.565 19.645 41.725 ;
        RECT 19.665 41.570 19.895 41.725 ;
        RECT 19.910 41.570 28.995 41.735 ;
        RECT 19.665 41.565 28.995 41.570 ;
        RECT 13.425 18.315 28.995 41.565 ;
        RECT 31.975 14.100 36.210 42.470 ;
      LAYER nwell ;
        RECT 36.470 42.380 39.630 46.535 ;
        RECT 36.435 36.455 39.625 40.415 ;
        RECT 36.435 30.005 39.625 33.965 ;
      LAYER pwell ;
        RECT 89.180 30.135 94.280 37.095 ;
      LAYER nwell ;
        RECT 36.435 23.555 39.625 27.515 ;
      LAYER pwell ;
        RECT 95.480 27.480 123.115 45.255 ;
        RECT 95.900 27.310 96.015 27.480 ;
        RECT 96.485 27.310 122.650 27.320 ;
      LAYER nwell ;
        RECT 36.515 14.170 39.690 21.035 ;
      LAYER li1 ;
        RECT 86.135 148.245 99.460 149.415 ;
        RECT 43.285 137.230 84.165 138.920 ;
        RECT 43.285 131.385 44.555 137.230 ;
        RECT 45.760 136.785 63.760 136.955 ;
        RECT 64.050 136.785 82.050 136.955 ;
        RECT 45.530 134.730 45.700 136.570 ;
        RECT 63.820 134.730 63.990 136.570 ;
        RECT 82.110 134.730 82.280 136.570 ;
        RECT 45.760 134.345 63.760 134.515 ;
        RECT 64.050 134.345 82.050 134.515 ;
        RECT 45.530 132.290 45.700 134.130 ;
        RECT 63.820 132.290 63.990 134.130 ;
        RECT 82.110 132.290 82.280 134.130 ;
        RECT 45.760 131.905 63.760 132.075 ;
        RECT 64.050 131.905 82.050 132.075 ;
        RECT 83.115 131.385 84.160 137.230 ;
        RECT 43.285 130.720 84.160 131.385 ;
        RECT 43.290 127.845 79.035 128.545 ;
        RECT 43.290 120.140 50.670 127.845 ;
        RECT 51.810 127.380 63.810 127.550 ;
        RECT 64.100 127.380 76.100 127.550 ;
        RECT 51.580 121.170 51.750 127.210 ;
        RECT 63.870 121.170 64.040 127.210 ;
        RECT 76.160 121.170 76.330 127.210 ;
        RECT 51.810 120.830 63.810 121.000 ;
        RECT 64.100 120.830 76.100 121.000 ;
        RECT 43.285 119.955 50.670 120.140 ;
        RECT 43.285 113.725 44.340 119.955 ;
        RECT 44.865 119.395 47.905 119.565 ;
        RECT 44.525 114.335 44.695 119.335 ;
        RECT 48.075 114.335 48.245 119.335 ;
        RECT 44.865 113.725 47.905 114.275 ;
        RECT 48.545 113.725 50.670 119.955 ;
        RECT 51.805 118.005 63.805 118.175 ;
        RECT 64.095 118.005 76.095 118.175 ;
        RECT 43.285 112.575 50.670 113.725 ;
        RECT 43.275 111.175 50.670 112.575 ;
        RECT 51.575 111.795 51.745 117.835 ;
        RECT 63.865 111.795 64.035 117.835 ;
        RECT 76.155 111.795 76.325 117.835 ;
        RECT 51.805 111.455 63.805 111.625 ;
        RECT 64.095 111.455 76.095 111.625 ;
        RECT 77.285 111.175 79.035 127.845 ;
        RECT 43.275 109.625 79.035 111.175 ;
        RECT 86.135 111.230 87.305 148.245 ;
        RECT 88.225 147.165 90.125 147.335 ;
        RECT 90.415 147.165 92.315 147.335 ;
        RECT 92.605 147.165 94.505 147.335 ;
        RECT 94.795 147.165 96.695 147.335 ;
        RECT 87.995 131.910 88.165 146.950 ;
        RECT 90.185 131.910 90.355 146.950 ;
        RECT 92.375 131.910 92.545 146.950 ;
        RECT 94.565 131.910 94.735 146.950 ;
        RECT 96.755 131.910 96.925 146.950 ;
        RECT 88.225 131.525 90.125 131.695 ;
        RECT 90.415 131.525 92.315 131.695 ;
        RECT 92.605 131.525 94.505 131.695 ;
        RECT 94.795 131.525 96.695 131.695 ;
        RECT 88.225 127.280 90.125 127.450 ;
        RECT 90.415 127.280 92.315 127.450 ;
        RECT 92.605 127.280 94.505 127.450 ;
        RECT 94.795 127.280 96.695 127.450 ;
        RECT 87.995 112.025 88.165 127.065 ;
        RECT 90.185 112.025 90.355 127.065 ;
        RECT 92.375 112.025 92.545 127.065 ;
        RECT 94.565 112.025 94.735 127.065 ;
        RECT 96.755 112.025 96.925 127.065 ;
        RECT 97.880 122.220 99.460 148.245 ;
        RECT 97.880 119.890 123.160 122.220 ;
        RECT 88.225 111.640 90.125 111.810 ;
        RECT 90.415 111.640 92.315 111.810 ;
        RECT 92.605 111.640 94.505 111.810 ;
        RECT 94.795 111.640 96.695 111.810 ;
        RECT 97.880 111.230 99.460 119.890 ;
        RECT 86.135 110.540 99.460 111.230 ;
        RECT 110.080 111.675 111.790 119.890 ;
        RECT 112.370 119.510 114.170 119.680 ;
        RECT 114.460 119.510 116.260 119.680 ;
        RECT 116.550 119.510 118.350 119.680 ;
        RECT 118.640 119.510 120.440 119.680 ;
        RECT 112.140 112.255 112.310 119.295 ;
        RECT 114.230 112.255 114.400 119.295 ;
        RECT 116.320 112.255 116.490 119.295 ;
        RECT 118.410 112.255 118.580 119.295 ;
        RECT 120.500 112.255 120.670 119.295 ;
        RECT 112.370 111.870 114.170 112.040 ;
        RECT 114.460 111.870 116.260 112.040 ;
        RECT 116.550 111.870 118.350 112.040 ;
        RECT 118.640 111.870 120.440 112.040 ;
        RECT 120.990 111.675 123.160 119.890 ;
        RECT 110.080 111.575 123.160 111.675 ;
        RECT 125.710 119.665 128.295 120.095 ;
        RECT 125.710 113.685 126.495 119.665 ;
        RECT 126.800 117.050 127.150 119.210 ;
        RECT 126.800 114.050 127.150 116.210 ;
        RECT 127.510 113.685 128.295 119.665 ;
        RECT 125.710 113.255 128.295 113.685 ;
        RECT 86.135 110.405 99.390 110.540 ;
        RECT 110.080 110.295 123.180 111.575 ;
        RECT 125.710 108.935 126.495 113.255 ;
        RECT 86.615 108.000 128.650 108.935 ;
        RECT 86.615 102.610 87.505 108.000 ;
        RECT 88.275 107.105 97.675 107.275 ;
        RECT 97.965 107.105 107.365 107.275 ;
        RECT 107.655 107.105 117.055 107.275 ;
        RECT 117.345 107.105 126.745 107.275 ;
        RECT 88.045 105.395 88.215 106.935 ;
        RECT 97.735 105.395 97.905 106.935 ;
        RECT 107.425 105.395 107.595 106.935 ;
        RECT 117.115 105.395 117.285 106.935 ;
        RECT 126.805 105.395 126.975 106.935 ;
        RECT 88.275 105.055 97.675 105.225 ;
        RECT 97.965 105.055 107.365 105.225 ;
        RECT 107.655 105.055 117.055 105.225 ;
        RECT 117.345 105.055 126.745 105.225 ;
        RECT 88.045 103.345 88.215 104.885 ;
        RECT 97.735 103.345 97.905 104.885 ;
        RECT 107.425 103.345 107.595 104.885 ;
        RECT 117.115 103.345 117.285 104.885 ;
        RECT 126.805 103.345 126.975 104.885 ;
        RECT 88.275 103.005 97.675 103.175 ;
        RECT 97.965 103.005 107.365 103.175 ;
        RECT 107.655 103.005 117.055 103.175 ;
        RECT 117.345 103.005 126.745 103.175 ;
        RECT 127.805 102.610 128.650 108.000 ;
        RECT 86.615 101.165 128.650 102.610 ;
        RECT 86.660 101.160 128.650 101.165 ;
        RECT 79.825 98.980 108.190 98.985 ;
        RECT 79.825 96.945 117.820 98.980 ;
        RECT 79.820 96.865 117.820 96.945 ;
        RECT 79.820 94.620 80.340 96.865 ;
        RECT 86.255 96.860 89.705 96.865 ;
        RECT 92.205 96.860 96.070 96.865 ;
        RECT 80.845 96.455 82.845 96.625 ;
        RECT 83.750 96.455 85.750 96.625 ;
        RECT 80.615 95.200 80.785 96.240 ;
        RECT 82.905 95.200 83.075 96.240 ;
        RECT 83.520 95.200 83.690 96.240 ;
        RECT 85.810 95.200 85.980 96.240 ;
        RECT 86.255 95.055 89.700 96.860 ;
        RECT 90.200 96.455 92.200 96.625 ;
        RECT 89.970 95.200 90.140 96.240 ;
        RECT 92.260 95.200 92.430 96.240 ;
        RECT 80.845 94.815 82.845 94.985 ;
        RECT 83.750 94.815 85.750 94.985 ;
        RECT 86.255 94.620 86.680 95.055 ;
        RECT 79.820 94.235 86.680 94.620 ;
        RECT 89.220 94.595 89.700 95.055 ;
        RECT 92.685 95.055 96.070 96.860 ;
        RECT 96.650 96.455 98.650 96.625 ;
        RECT 96.420 95.200 96.590 96.240 ;
        RECT 98.710 95.200 98.880 96.240 ;
        RECT 90.200 94.815 92.200 94.985 ;
        RECT 92.685 94.595 93.140 95.055 ;
        RECT 79.820 94.225 86.670 94.235 ;
        RECT 89.220 94.180 93.140 94.595 ;
        RECT 95.670 94.605 96.070 95.055 ;
        RECT 99.175 95.115 102.565 96.865 ;
        RECT 105.625 96.825 117.820 96.865 ;
        RECT 103.100 96.455 105.100 96.625 ;
        RECT 102.870 95.200 103.040 96.240 ;
        RECT 105.160 95.200 105.330 96.240 ;
        RECT 96.650 94.815 98.650 94.985 ;
        RECT 99.175 94.605 99.600 95.115 ;
        RECT 95.670 94.225 99.620 94.605 ;
        RECT 102.175 94.535 102.565 95.115 ;
        RECT 103.100 94.815 105.100 94.985 ;
        RECT 105.625 94.535 106.015 96.825 ;
        RECT 102.170 94.205 106.015 94.535 ;
        RECT 107.730 94.590 107.975 96.825 ;
        RECT 111.450 96.815 117.820 96.825 ;
        RECT 111.450 96.810 116.390 96.815 ;
        RECT 116.620 96.810 117.820 96.815 ;
        RECT 108.540 96.455 109.540 96.625 ;
        RECT 109.830 96.455 110.830 96.625 ;
        RECT 108.310 95.200 108.480 96.240 ;
        RECT 109.600 95.200 109.770 96.240 ;
        RECT 110.890 95.200 111.060 96.240 ;
        RECT 112.165 95.955 114.165 96.125 ;
        RECT 114.455 95.955 116.455 96.125 ;
        RECT 111.935 95.200 112.105 95.740 ;
        RECT 114.225 95.200 114.395 95.740 ;
        RECT 116.515 95.200 116.685 95.740 ;
        RECT 108.540 94.815 109.540 94.985 ;
        RECT 109.830 94.815 110.830 94.985 ;
        RECT 112.165 94.815 114.165 94.985 ;
        RECT 114.455 94.815 116.455 94.985 ;
        RECT 117.175 94.590 117.435 96.810 ;
        RECT 107.730 94.350 117.435 94.590 ;
        RECT 102.170 94.195 106.005 94.205 ;
        RECT 79.870 93.160 107.980 93.855 ;
        RECT 79.870 90.685 80.485 93.160 ;
        RECT 81.170 92.475 82.170 92.645 ;
        RECT 82.460 92.475 83.460 92.645 ;
        RECT 83.750 92.475 84.750 92.645 ;
        RECT 85.040 92.475 86.040 92.645 ;
        RECT 86.330 92.475 87.330 92.645 ;
        RECT 87.620 92.475 88.620 92.645 ;
        RECT 88.910 92.475 89.910 92.645 ;
        RECT 90.200 92.475 91.200 92.645 ;
        RECT 91.490 92.475 92.490 92.645 ;
        RECT 92.780 92.475 93.780 92.645 ;
        RECT 94.070 92.475 95.070 92.645 ;
        RECT 95.360 92.475 96.360 92.645 ;
        RECT 96.650 92.475 97.650 92.645 ;
        RECT 97.940 92.475 98.940 92.645 ;
        RECT 99.230 92.475 100.230 92.645 ;
        RECT 100.520 92.475 101.520 92.645 ;
        RECT 101.810 92.475 102.810 92.645 ;
        RECT 103.100 92.475 104.100 92.645 ;
        RECT 104.390 92.475 105.390 92.645 ;
        RECT 105.680 92.475 106.680 92.645 ;
        RECT 80.940 91.265 81.110 92.305 ;
        RECT 82.230 91.265 82.400 92.305 ;
        RECT 83.520 91.265 83.690 92.305 ;
        RECT 84.810 91.265 84.980 92.305 ;
        RECT 86.100 91.265 86.270 92.305 ;
        RECT 87.390 91.265 87.560 92.305 ;
        RECT 88.680 91.265 88.850 92.305 ;
        RECT 89.970 91.265 90.140 92.305 ;
        RECT 91.260 91.265 91.430 92.305 ;
        RECT 92.550 91.265 92.720 92.305 ;
        RECT 93.840 91.265 94.010 92.305 ;
        RECT 95.130 91.265 95.300 92.305 ;
        RECT 96.420 91.265 96.590 92.305 ;
        RECT 97.710 91.265 97.880 92.305 ;
        RECT 99.000 91.265 99.170 92.305 ;
        RECT 100.290 91.265 100.460 92.305 ;
        RECT 101.580 91.265 101.750 92.305 ;
        RECT 102.870 91.265 103.040 92.305 ;
        RECT 104.160 91.265 104.330 92.305 ;
        RECT 105.450 91.265 105.620 92.305 ;
        RECT 106.740 91.265 106.910 92.305 ;
        RECT 81.170 90.925 82.170 91.095 ;
        RECT 82.460 90.925 83.460 91.095 ;
        RECT 83.750 90.925 84.750 91.095 ;
        RECT 85.040 90.925 86.040 91.095 ;
        RECT 86.330 90.925 87.330 91.095 ;
        RECT 87.620 90.925 88.620 91.095 ;
        RECT 88.910 90.925 89.910 91.095 ;
        RECT 90.200 90.925 91.200 91.095 ;
        RECT 91.490 90.925 92.490 91.095 ;
        RECT 92.780 90.925 93.780 91.095 ;
        RECT 94.070 90.925 95.070 91.095 ;
        RECT 95.360 90.925 96.360 91.095 ;
        RECT 96.650 90.925 97.650 91.095 ;
        RECT 97.940 90.925 98.940 91.095 ;
        RECT 99.230 90.925 100.230 91.095 ;
        RECT 100.520 90.925 101.520 91.095 ;
        RECT 101.810 90.925 102.810 91.095 ;
        RECT 103.100 90.925 104.100 91.095 ;
        RECT 104.390 90.925 105.390 91.095 ;
        RECT 105.680 90.925 106.680 91.095 ;
        RECT 107.365 90.685 107.980 93.160 ;
        RECT 79.870 89.460 107.980 90.685 ;
        RECT 110.855 92.310 117.295 93.485 ;
        RECT 79.870 89.405 108.005 89.460 ;
        RECT 84.115 87.075 108.005 89.405 ;
        RECT 110.855 88.220 112.030 92.310 ;
        RECT 112.340 88.530 115.810 92.000 ;
        RECT 116.120 88.220 117.295 92.310 ;
        RECT 110.855 87.075 117.295 88.220 ;
        RECT 84.115 87.045 117.295 87.075 ;
        RECT 84.115 86.640 117.290 87.045 ;
        RECT 84.130 86.615 117.290 86.640 ;
        RECT 84.130 85.610 117.285 86.615 ;
        RECT 84.130 85.575 116.025 85.610 ;
        RECT 84.130 72.545 84.710 85.575 ;
        RECT 85.195 84.790 86.195 84.960 ;
        RECT 86.485 84.790 87.485 84.960 ;
        RECT 87.775 84.790 88.775 84.960 ;
        RECT 89.065 84.790 90.065 84.960 ;
        RECT 90.355 84.790 91.355 84.960 ;
        RECT 91.645 84.790 92.645 84.960 ;
        RECT 92.935 84.790 93.935 84.960 ;
        RECT 94.225 84.790 95.225 84.960 ;
        RECT 95.515 84.790 96.515 84.960 ;
        RECT 96.805 84.790 97.805 84.960 ;
        RECT 98.095 84.790 99.095 84.960 ;
        RECT 99.385 84.790 100.385 84.960 ;
        RECT 100.675 84.790 101.675 84.960 ;
        RECT 101.965 84.790 102.965 84.960 ;
        RECT 103.255 84.790 104.255 84.960 ;
        RECT 104.545 84.790 105.545 84.960 ;
        RECT 105.835 84.790 106.835 84.960 ;
        RECT 107.125 84.790 108.125 84.960 ;
        RECT 108.415 84.790 109.415 84.960 ;
        RECT 109.705 84.790 110.705 84.960 ;
        RECT 110.995 84.790 111.995 84.960 ;
        RECT 112.285 84.790 113.285 84.960 ;
        RECT 113.575 84.790 114.575 84.960 ;
        RECT 114.865 84.790 115.865 84.960 ;
        RECT 84.965 80.580 85.135 84.620 ;
        RECT 86.255 80.580 86.425 84.620 ;
        RECT 87.545 80.580 87.715 84.620 ;
        RECT 88.835 80.580 89.005 84.620 ;
        RECT 90.125 80.580 90.295 84.620 ;
        RECT 91.415 80.580 91.585 84.620 ;
        RECT 92.705 80.580 92.875 84.620 ;
        RECT 93.995 80.580 94.165 84.620 ;
        RECT 95.285 80.580 95.455 84.620 ;
        RECT 96.575 80.580 96.745 84.620 ;
        RECT 97.865 80.580 98.035 84.620 ;
        RECT 99.155 80.580 99.325 84.620 ;
        RECT 100.445 80.580 100.615 84.620 ;
        RECT 101.735 80.580 101.905 84.620 ;
        RECT 103.025 80.580 103.195 84.620 ;
        RECT 104.315 80.580 104.485 84.620 ;
        RECT 105.605 80.580 105.775 84.620 ;
        RECT 106.895 80.580 107.065 84.620 ;
        RECT 108.185 80.580 108.355 84.620 ;
        RECT 109.475 80.580 109.645 84.620 ;
        RECT 110.765 80.580 110.935 84.620 ;
        RECT 112.055 80.580 112.225 84.620 ;
        RECT 113.345 80.580 113.515 84.620 ;
        RECT 114.635 80.580 114.805 84.620 ;
        RECT 115.925 80.580 116.095 84.620 ;
        RECT 85.195 80.240 86.195 80.410 ;
        RECT 86.485 80.240 87.485 80.410 ;
        RECT 87.775 80.240 88.775 80.410 ;
        RECT 89.065 80.240 90.065 80.410 ;
        RECT 90.355 80.240 91.355 80.410 ;
        RECT 91.645 80.240 92.645 80.410 ;
        RECT 92.935 80.240 93.935 80.410 ;
        RECT 94.225 80.240 95.225 80.410 ;
        RECT 95.515 80.240 96.515 80.410 ;
        RECT 96.805 80.240 97.805 80.410 ;
        RECT 98.095 80.240 99.095 80.410 ;
        RECT 99.385 80.240 100.385 80.410 ;
        RECT 100.675 80.240 101.675 80.410 ;
        RECT 101.965 80.240 102.965 80.410 ;
        RECT 103.255 80.240 104.255 80.410 ;
        RECT 104.545 80.240 105.545 80.410 ;
        RECT 105.835 80.240 106.835 80.410 ;
        RECT 107.125 80.240 108.125 80.410 ;
        RECT 108.415 80.240 109.415 80.410 ;
        RECT 109.705 80.240 110.705 80.410 ;
        RECT 110.995 80.240 111.995 80.410 ;
        RECT 112.285 80.240 113.285 80.410 ;
        RECT 113.575 80.240 114.575 80.410 ;
        RECT 114.865 80.240 115.865 80.410 ;
        RECT 85.195 77.385 86.195 77.555 ;
        RECT 86.485 77.385 87.485 77.555 ;
        RECT 87.775 77.385 88.775 77.555 ;
        RECT 89.065 77.385 90.065 77.555 ;
        RECT 90.355 77.385 91.355 77.555 ;
        RECT 91.645 77.385 92.645 77.555 ;
        RECT 92.935 77.385 93.935 77.555 ;
        RECT 94.225 77.385 95.225 77.555 ;
        RECT 95.515 77.385 96.515 77.555 ;
        RECT 96.805 77.385 97.805 77.555 ;
        RECT 98.095 77.385 99.095 77.555 ;
        RECT 99.385 77.385 100.385 77.555 ;
        RECT 100.675 77.385 101.675 77.555 ;
        RECT 101.965 77.385 102.965 77.555 ;
        RECT 103.255 77.385 104.255 77.555 ;
        RECT 104.545 77.385 105.545 77.555 ;
        RECT 105.835 77.385 106.835 77.555 ;
        RECT 107.125 77.385 108.125 77.555 ;
        RECT 108.415 77.385 109.415 77.555 ;
        RECT 109.705 77.385 110.705 77.555 ;
        RECT 110.995 77.385 111.995 77.555 ;
        RECT 112.285 77.385 113.285 77.555 ;
        RECT 113.575 77.385 114.575 77.555 ;
        RECT 114.865 77.385 115.865 77.555 ;
        RECT 84.965 73.175 85.135 77.215 ;
        RECT 86.255 73.175 86.425 77.215 ;
        RECT 87.545 73.175 87.715 77.215 ;
        RECT 88.835 73.175 89.005 77.215 ;
        RECT 90.125 73.175 90.295 77.215 ;
        RECT 91.415 73.175 91.585 77.215 ;
        RECT 92.705 73.175 92.875 77.215 ;
        RECT 93.995 73.175 94.165 77.215 ;
        RECT 95.285 73.175 95.455 77.215 ;
        RECT 96.575 73.175 96.745 77.215 ;
        RECT 97.865 73.175 98.035 77.215 ;
        RECT 99.155 73.175 99.325 77.215 ;
        RECT 100.445 73.175 100.615 77.215 ;
        RECT 101.735 73.175 101.905 77.215 ;
        RECT 103.025 73.175 103.195 77.215 ;
        RECT 104.315 73.175 104.485 77.215 ;
        RECT 105.605 73.175 105.775 77.215 ;
        RECT 106.895 73.175 107.065 77.215 ;
        RECT 108.185 73.175 108.355 77.215 ;
        RECT 109.475 73.175 109.645 77.215 ;
        RECT 110.765 73.175 110.935 77.215 ;
        RECT 112.055 73.175 112.225 77.215 ;
        RECT 113.345 73.175 113.515 77.215 ;
        RECT 114.635 73.175 114.805 77.215 ;
        RECT 115.925 73.175 116.095 77.215 ;
        RECT 85.195 72.835 86.195 73.005 ;
        RECT 86.485 72.835 87.485 73.005 ;
        RECT 87.775 72.835 88.775 73.005 ;
        RECT 89.065 72.835 90.065 73.005 ;
        RECT 90.355 72.835 91.355 73.005 ;
        RECT 91.645 72.835 92.645 73.005 ;
        RECT 92.935 72.835 93.935 73.005 ;
        RECT 94.225 72.835 95.225 73.005 ;
        RECT 95.515 72.835 96.515 73.005 ;
        RECT 96.805 72.835 97.805 73.005 ;
        RECT 98.095 72.835 99.095 73.005 ;
        RECT 99.385 72.835 100.385 73.005 ;
        RECT 100.675 72.835 101.675 73.005 ;
        RECT 101.965 72.835 102.965 73.005 ;
        RECT 103.255 72.835 104.255 73.005 ;
        RECT 104.545 72.835 105.545 73.005 ;
        RECT 105.835 72.835 106.835 73.005 ;
        RECT 107.125 72.835 108.125 73.005 ;
        RECT 108.415 72.835 109.415 73.005 ;
        RECT 109.705 72.835 110.705 73.005 ;
        RECT 110.995 72.835 111.995 73.005 ;
        RECT 112.285 72.835 113.285 73.005 ;
        RECT 113.575 72.835 114.575 73.005 ;
        RECT 114.865 72.835 115.865 73.005 ;
        RECT 116.825 72.545 117.285 85.610 ;
        RECT 84.130 70.740 117.720 72.545 ;
        RECT 88.630 54.010 129.510 55.700 ;
        RECT 13.050 52.115 14.855 52.550 ;
        RECT 39.120 52.265 41.290 52.650 ;
        RECT 29.355 52.120 35.795 52.125 ;
        RECT 28.925 52.115 35.795 52.120 ;
        RECT 13.050 51.655 35.795 52.115 ;
        RECT 13.050 19.540 14.855 51.655 ;
        RECT 27.920 50.950 35.795 51.655 ;
        RECT 15.485 50.755 19.525 50.925 ;
        RECT 22.890 50.755 26.930 50.925 ;
        RECT 27.920 50.855 30.530 50.950 ;
        RECT 15.145 49.695 15.315 50.695 ;
        RECT 19.695 49.695 19.865 50.695 ;
        RECT 22.550 49.695 22.720 50.695 ;
        RECT 27.100 49.695 27.270 50.695 ;
        RECT 15.485 49.465 19.525 49.635 ;
        RECT 22.890 49.465 26.930 49.635 ;
        RECT 15.145 48.405 15.315 49.405 ;
        RECT 19.695 48.405 19.865 49.405 ;
        RECT 22.550 48.405 22.720 49.405 ;
        RECT 27.100 48.405 27.270 49.405 ;
        RECT 15.485 48.175 19.525 48.345 ;
        RECT 22.890 48.175 26.930 48.345 ;
        RECT 15.145 47.115 15.315 48.115 ;
        RECT 19.695 47.115 19.865 48.115 ;
        RECT 22.550 47.115 22.720 48.115 ;
        RECT 27.100 47.115 27.270 48.115 ;
        RECT 15.485 46.885 19.525 47.055 ;
        RECT 22.890 46.885 26.930 47.055 ;
        RECT 27.885 46.860 30.530 50.855 ;
        RECT 30.840 47.170 34.310 50.640 ;
        RECT 34.620 46.860 35.795 50.950 ;
        RECT 15.145 45.825 15.315 46.825 ;
        RECT 19.695 45.825 19.865 46.825 ;
        RECT 22.550 45.825 22.720 46.825 ;
        RECT 27.100 45.825 27.270 46.825 ;
        RECT 15.485 45.595 19.525 45.765 ;
        RECT 22.890 45.595 26.930 45.765 ;
        RECT 27.885 45.685 35.795 46.860 ;
        RECT 36.660 52.005 41.290 52.265 ;
        RECT 15.145 44.535 15.315 45.535 ;
        RECT 19.695 44.535 19.865 45.535 ;
        RECT 22.550 44.535 22.720 45.535 ;
        RECT 27.100 44.535 27.270 45.535 ;
        RECT 15.485 44.305 19.525 44.475 ;
        RECT 22.890 44.305 26.930 44.475 ;
        RECT 15.145 43.245 15.315 44.245 ;
        RECT 19.695 43.245 19.865 44.245 ;
        RECT 22.550 43.245 22.720 44.245 ;
        RECT 27.100 43.245 27.270 44.245 ;
        RECT 15.485 43.015 19.525 43.185 ;
        RECT 22.890 43.015 26.930 43.185 ;
        RECT 15.145 41.955 15.315 42.955 ;
        RECT 19.695 41.955 19.865 42.955 ;
        RECT 22.550 41.955 22.720 42.955 ;
        RECT 27.100 41.955 27.270 42.955 ;
        RECT 27.885 42.320 29.385 45.685 ;
        RECT 36.660 42.805 36.900 52.005 ;
        RECT 37.510 51.345 38.050 51.515 ;
        RECT 39.120 51.450 41.290 52.005 ;
        RECT 37.125 49.285 37.295 51.285 ;
        RECT 38.265 49.285 38.435 51.285 ;
        RECT 39.125 51.220 41.290 51.450 ;
        RECT 37.510 49.055 38.050 49.225 ;
        RECT 37.125 46.995 37.295 48.995 ;
        RECT 38.265 46.995 38.435 48.995 ;
        RECT 37.510 46.765 38.050 46.935 ;
        RECT 39.120 46.280 41.290 51.220 ;
        RECT 88.630 48.165 89.900 54.010 ;
        RECT 91.105 53.565 109.105 53.735 ;
        RECT 109.395 53.565 127.395 53.735 ;
        RECT 90.875 51.510 91.045 53.350 ;
        RECT 109.165 51.510 109.335 53.350 ;
        RECT 127.455 51.510 127.625 53.350 ;
        RECT 91.105 51.125 109.105 51.295 ;
        RECT 109.395 51.125 127.395 51.295 ;
        RECT 90.875 49.070 91.045 50.910 ;
        RECT 109.165 49.070 109.335 50.910 ;
        RECT 127.455 49.070 127.625 50.910 ;
        RECT 91.105 48.685 109.105 48.855 ;
        RECT 109.395 48.685 127.395 48.855 ;
        RECT 128.460 48.165 129.505 54.010 ;
        RECT 88.630 47.500 129.505 48.165 ;
        RECT 37.510 45.720 38.550 45.890 ;
        RECT 37.125 44.660 37.295 45.660 ;
        RECT 38.765 44.660 38.935 45.660 ;
        RECT 37.510 44.430 38.550 44.600 ;
        RECT 37.125 43.370 37.295 44.370 ;
        RECT 38.765 43.370 38.935 44.370 ;
        RECT 37.510 43.140 38.550 43.310 ;
        RECT 39.135 42.805 41.290 46.280 ;
        RECT 36.660 42.560 41.290 42.805 ;
        RECT 39.135 42.385 41.290 42.560 ;
        RECT 88.635 44.625 124.380 45.325 ;
        RECT 27.885 42.315 31.760 42.320 ;
        RECT 15.485 41.725 19.525 41.895 ;
        RECT 22.890 41.725 26.930 41.895 ;
        RECT 27.885 41.700 36.165 42.315 ;
        RECT 15.145 40.665 15.315 41.665 ;
        RECT 19.695 40.665 19.865 41.665 ;
        RECT 22.550 40.665 22.720 41.665 ;
        RECT 27.100 40.665 27.270 41.665 ;
        RECT 15.485 40.435 19.525 40.605 ;
        RECT 22.890 40.435 26.930 40.605 ;
        RECT 15.145 39.375 15.315 40.375 ;
        RECT 19.695 39.375 19.865 40.375 ;
        RECT 22.550 39.375 22.720 40.375 ;
        RECT 27.100 39.375 27.270 40.375 ;
        RECT 15.485 39.145 19.525 39.315 ;
        RECT 22.890 39.145 26.930 39.315 ;
        RECT 15.145 38.085 15.315 39.085 ;
        RECT 19.695 38.085 19.865 39.085 ;
        RECT 22.550 38.085 22.720 39.085 ;
        RECT 27.100 38.085 27.270 39.085 ;
        RECT 15.485 37.855 19.525 38.025 ;
        RECT 22.890 37.855 26.930 38.025 ;
        RECT 15.145 36.795 15.315 37.795 ;
        RECT 19.695 36.795 19.865 37.795 ;
        RECT 22.550 36.795 22.720 37.795 ;
        RECT 27.100 36.795 27.270 37.795 ;
        RECT 15.485 36.565 19.525 36.735 ;
        RECT 22.890 36.565 26.930 36.735 ;
        RECT 15.145 35.505 15.315 36.505 ;
        RECT 19.695 35.505 19.865 36.505 ;
        RECT 22.550 35.505 22.720 36.505 ;
        RECT 27.100 35.505 27.270 36.505 ;
        RECT 15.485 35.275 19.525 35.445 ;
        RECT 22.890 35.275 26.930 35.445 ;
        RECT 15.145 34.215 15.315 35.215 ;
        RECT 19.695 34.215 19.865 35.215 ;
        RECT 22.550 34.215 22.720 35.215 ;
        RECT 27.100 34.215 27.270 35.215 ;
        RECT 15.485 33.985 19.525 34.155 ;
        RECT 22.890 33.985 26.930 34.155 ;
        RECT 15.145 32.925 15.315 33.925 ;
        RECT 19.695 32.925 19.865 33.925 ;
        RECT 22.550 32.925 22.720 33.925 ;
        RECT 27.100 32.925 27.270 33.925 ;
        RECT 15.485 32.695 19.525 32.865 ;
        RECT 22.890 32.695 26.930 32.865 ;
        RECT 15.145 31.635 15.315 32.635 ;
        RECT 19.695 31.635 19.865 32.635 ;
        RECT 22.550 31.635 22.720 32.635 ;
        RECT 27.100 31.635 27.270 32.635 ;
        RECT 15.485 31.405 19.525 31.575 ;
        RECT 22.890 31.405 26.930 31.575 ;
        RECT 15.145 30.345 15.315 31.345 ;
        RECT 19.695 30.345 19.865 31.345 ;
        RECT 22.550 30.345 22.720 31.345 ;
        RECT 27.100 30.345 27.270 31.345 ;
        RECT 15.485 30.115 19.525 30.285 ;
        RECT 22.890 30.115 26.930 30.285 ;
        RECT 15.145 29.055 15.315 30.055 ;
        RECT 19.695 29.055 19.865 30.055 ;
        RECT 22.550 29.055 22.720 30.055 ;
        RECT 27.100 29.055 27.270 30.055 ;
        RECT 15.485 28.825 19.525 28.995 ;
        RECT 22.890 28.825 26.930 28.995 ;
        RECT 15.145 27.765 15.315 28.765 ;
        RECT 19.695 27.765 19.865 28.765 ;
        RECT 22.550 27.765 22.720 28.765 ;
        RECT 27.100 27.765 27.270 28.765 ;
        RECT 15.485 27.535 19.525 27.705 ;
        RECT 22.890 27.535 26.930 27.705 ;
        RECT 15.145 26.475 15.315 27.475 ;
        RECT 19.695 26.475 19.865 27.475 ;
        RECT 22.550 26.475 22.720 27.475 ;
        RECT 27.100 26.475 27.270 27.475 ;
        RECT 15.485 26.245 19.525 26.415 ;
        RECT 22.890 26.245 26.930 26.415 ;
        RECT 15.145 25.185 15.315 26.185 ;
        RECT 19.695 25.185 19.865 26.185 ;
        RECT 22.550 25.185 22.720 26.185 ;
        RECT 27.100 25.185 27.270 26.185 ;
        RECT 15.485 24.955 19.525 25.125 ;
        RECT 22.890 24.955 26.930 25.125 ;
        RECT 15.145 23.895 15.315 24.895 ;
        RECT 19.695 23.895 19.865 24.895 ;
        RECT 22.550 23.895 22.720 24.895 ;
        RECT 27.100 23.895 27.270 24.895 ;
        RECT 15.485 23.665 19.525 23.835 ;
        RECT 22.890 23.665 26.930 23.835 ;
        RECT 15.145 22.605 15.315 23.605 ;
        RECT 19.695 22.605 19.865 23.605 ;
        RECT 22.550 22.605 22.720 23.605 ;
        RECT 27.100 22.605 27.270 23.605 ;
        RECT 15.485 22.375 19.525 22.545 ;
        RECT 22.890 22.375 26.930 22.545 ;
        RECT 15.145 21.315 15.315 22.315 ;
        RECT 19.695 21.315 19.865 22.315 ;
        RECT 22.550 21.315 22.720 22.315 ;
        RECT 27.100 21.315 27.270 22.315 ;
        RECT 15.485 21.085 19.525 21.255 ;
        RECT 22.890 21.085 26.930 21.255 ;
        RECT 15.145 20.025 15.315 21.025 ;
        RECT 19.695 20.025 19.865 21.025 ;
        RECT 22.550 20.025 22.720 21.025 ;
        RECT 27.100 20.025 27.270 21.025 ;
        RECT 15.485 19.795 19.525 19.965 ;
        RECT 22.890 19.795 26.930 19.965 ;
        RECT 27.885 19.540 32.995 41.700 ;
        RECT 33.575 41.075 34.615 41.245 ;
        RECT 33.235 40.015 33.405 41.015 ;
        RECT 34.785 40.015 34.955 41.015 ;
        RECT 33.575 39.785 34.615 39.955 ;
        RECT 33.235 38.725 33.405 39.725 ;
        RECT 34.785 38.725 34.955 39.725 ;
        RECT 33.575 38.495 34.615 38.665 ;
        RECT 33.235 37.435 33.405 38.435 ;
        RECT 34.785 37.435 34.955 38.435 ;
        RECT 33.575 37.205 34.615 37.375 ;
        RECT 33.235 36.145 33.405 37.145 ;
        RECT 34.785 36.145 34.955 37.145 ;
        RECT 33.575 35.915 34.615 36.085 ;
        RECT 33.235 34.855 33.405 35.855 ;
        RECT 34.785 34.855 34.955 35.855 ;
        RECT 33.575 34.625 34.615 34.795 ;
        RECT 33.235 33.565 33.405 34.565 ;
        RECT 34.785 33.565 34.955 34.565 ;
        RECT 33.575 33.335 34.615 33.505 ;
        RECT 33.235 32.275 33.405 33.275 ;
        RECT 34.785 32.275 34.955 33.275 ;
        RECT 33.575 32.045 34.615 32.215 ;
        RECT 33.235 30.985 33.405 31.985 ;
        RECT 34.785 30.985 34.955 31.985 ;
        RECT 33.575 30.755 34.615 30.925 ;
        RECT 33.235 29.695 33.405 30.695 ;
        RECT 34.785 29.695 34.955 30.695 ;
        RECT 33.575 29.465 34.615 29.635 ;
        RECT 33.235 28.405 33.405 29.405 ;
        RECT 34.785 28.405 34.955 29.405 ;
        RECT 33.575 28.175 34.615 28.345 ;
        RECT 33.235 27.115 33.405 28.115 ;
        RECT 34.785 27.115 34.955 28.115 ;
        RECT 33.575 26.885 34.615 27.055 ;
        RECT 33.235 25.825 33.405 26.825 ;
        RECT 34.785 25.825 34.955 26.825 ;
        RECT 33.575 25.595 34.615 25.765 ;
        RECT 33.235 24.535 33.405 25.535 ;
        RECT 34.785 24.535 34.955 25.535 ;
        RECT 33.575 24.305 34.615 24.475 ;
        RECT 33.235 23.245 33.405 24.245 ;
        RECT 34.785 23.245 34.955 24.245 ;
        RECT 33.575 23.015 34.615 23.185 ;
        RECT 33.235 21.955 33.405 22.955 ;
        RECT 34.785 21.955 34.955 22.955 ;
        RECT 33.575 21.725 34.615 21.895 ;
        RECT 33.235 20.665 33.405 21.665 ;
        RECT 34.785 20.665 34.955 21.665 ;
        RECT 33.575 20.435 34.615 20.605 ;
        RECT 13.050 18.960 32.995 19.540 ;
        RECT 33.235 19.375 33.405 20.375 ;
        RECT 34.785 19.375 34.955 20.375 ;
        RECT 33.575 19.145 34.615 19.315 ;
        RECT 31.715 14.820 32.995 18.960 ;
        RECT 33.235 18.085 33.405 19.085 ;
        RECT 34.785 18.085 34.955 19.085 ;
        RECT 33.575 17.855 34.615 18.025 ;
        RECT 33.235 16.795 33.405 17.795 ;
        RECT 34.785 16.795 34.955 17.795 ;
        RECT 33.575 16.565 34.615 16.735 ;
        RECT 33.235 15.505 33.405 16.505 ;
        RECT 34.785 15.505 34.955 16.505 ;
        RECT 33.575 15.275 34.615 15.445 ;
        RECT 35.470 14.820 36.165 41.700 ;
        RECT 36.515 40.340 40.800 40.350 ;
        RECT 36.505 39.960 40.800 40.340 ;
        RECT 36.505 36.900 36.845 39.960 ;
        RECT 37.510 39.495 38.550 39.665 ;
        RECT 37.125 37.435 37.295 39.435 ;
        RECT 38.765 37.435 38.935 39.435 ;
        RECT 37.510 37.205 38.550 37.375 ;
        RECT 39.175 36.900 40.800 39.960 ;
        RECT 88.635 36.920 96.015 44.625 ;
        RECT 97.155 44.160 109.155 44.330 ;
        RECT 109.445 44.160 121.445 44.330 ;
        RECT 96.925 37.950 97.095 43.990 ;
        RECT 109.215 37.950 109.385 43.990 ;
        RECT 121.505 37.950 121.675 43.990 ;
        RECT 97.155 37.610 109.155 37.780 ;
        RECT 109.445 37.610 121.445 37.780 ;
        RECT 36.505 36.510 40.800 36.900 ;
        RECT 36.505 36.505 36.845 36.510 ;
        RECT 36.535 33.935 36.915 33.955 ;
        RECT 37.425 33.935 40.800 36.510 ;
        RECT 36.535 33.510 40.800 33.935 ;
        RECT 36.535 30.405 36.915 33.510 ;
        RECT 37.510 33.045 38.550 33.215 ;
        RECT 37.125 30.985 37.295 32.985 ;
        RECT 38.765 30.985 38.935 32.985 ;
        RECT 37.510 30.755 38.550 30.925 ;
        RECT 39.175 30.405 40.800 33.510 ;
        RECT 36.535 30.005 40.800 30.405 ;
        RECT 37.365 27.475 40.800 30.005 ;
        RECT 88.630 36.735 96.015 36.920 ;
        RECT 88.630 30.505 89.685 36.735 ;
        RECT 90.210 36.175 93.250 36.345 ;
        RECT 89.870 31.115 90.040 36.115 ;
        RECT 93.420 31.115 93.590 36.115 ;
        RECT 90.210 30.505 93.250 31.055 ;
        RECT 93.890 30.505 96.015 36.735 ;
        RECT 97.150 34.785 109.150 34.955 ;
        RECT 109.440 34.785 121.440 34.955 ;
        RECT 88.630 29.355 96.015 30.505 ;
        RECT 36.490 27.020 40.800 27.475 ;
        RECT 36.490 24.035 36.905 27.020 ;
        RECT 37.510 26.595 38.550 26.765 ;
        RECT 39.170 26.540 40.800 27.020 ;
        RECT 37.125 24.535 37.295 26.535 ;
        RECT 38.765 24.535 38.935 26.535 ;
        RECT 37.510 24.305 38.550 24.475 ;
        RECT 39.175 24.040 40.800 26.540 ;
        RECT 88.620 27.955 96.015 29.355 ;
        RECT 96.920 28.575 97.090 34.615 ;
        RECT 109.210 28.575 109.380 34.615 ;
        RECT 121.500 28.575 121.670 34.615 ;
        RECT 97.150 28.235 109.150 28.405 ;
        RECT 109.440 28.235 121.440 28.405 ;
        RECT 122.630 27.955 124.380 44.625 ;
        RECT 88.620 26.405 124.380 27.955 ;
        RECT 39.170 24.035 40.800 24.040 ;
        RECT 36.490 23.555 40.800 24.035 ;
        RECT 37.365 21.370 40.800 23.555 ;
        RECT 37.365 21.015 40.805 21.370 ;
        RECT 36.545 21.005 40.805 21.015 ;
        RECT 31.715 14.205 36.165 14.820 ;
        RECT 36.535 20.590 40.805 21.005 ;
        RECT 36.535 14.675 36.930 20.590 ;
        RECT 37.510 20.145 38.550 20.315 ;
        RECT 37.125 18.085 37.295 20.085 ;
        RECT 38.765 18.085 38.935 20.085 ;
        RECT 37.510 17.855 38.550 18.025 ;
        RECT 37.510 17.240 38.550 17.410 ;
        RECT 37.125 15.180 37.295 17.180 ;
        RECT 38.765 15.180 38.935 17.180 ;
        RECT 37.510 14.950 38.550 15.120 ;
        RECT 39.175 14.675 40.805 20.590 ;
        RECT 36.535 14.160 40.805 14.675 ;
        RECT 36.535 14.155 39.255 14.160 ;
      LAYER met1 ;
        RECT 86.245 148.305 99.325 149.380 ;
        RECT 44.145 138.265 83.255 138.770 ;
        RECT 44.795 136.755 82.030 136.985 ;
        RECT 44.795 134.745 45.795 136.755 ;
        RECT 44.795 129.590 45.225 134.745 ;
        RECT 46.680 134.545 62.875 136.755 ;
        RECT 63.790 136.490 64.020 136.550 ;
        RECT 63.720 134.810 64.090 136.490 ;
        RECT 63.790 134.750 64.020 134.810 ;
        RECT 64.990 134.545 81.185 136.755 ;
        RECT 82.010 134.755 83.020 136.555 ;
        RECT 82.080 134.750 82.310 134.755 ;
        RECT 45.780 134.315 63.740 134.545 ;
        RECT 64.070 134.315 82.030 134.545 ;
        RECT 45.365 132.305 45.795 134.110 ;
        RECT 46.680 132.105 62.875 134.315 ;
        RECT 63.790 134.050 64.020 134.110 ;
        RECT 63.720 132.370 64.090 134.050 ;
        RECT 63.790 132.310 64.020 132.370 ;
        RECT 64.990 132.105 81.185 134.315 ;
        RECT 82.020 132.105 82.450 134.110 ;
        RECT 45.780 131.875 82.450 132.105 ;
        RECT 82.590 130.515 83.020 134.755 ;
        RECT 86.255 131.295 87.180 148.305 ;
        RECT 88.245 147.135 90.105 147.365 ;
        RECT 90.435 147.135 92.295 147.365 ;
        RECT 92.625 147.135 94.485 147.365 ;
        RECT 94.815 147.135 96.675 147.365 ;
        RECT 87.965 136.990 88.195 146.930 ;
        RECT 87.865 131.990 88.285 136.990 ;
        RECT 87.965 131.930 88.195 131.990 ;
        RECT 88.605 131.740 89.630 147.135 ;
        RECT 90.155 146.870 90.385 146.930 ;
        RECT 90.040 143.870 90.500 146.870 ;
        RECT 90.155 131.930 90.385 143.870 ;
        RECT 90.870 131.740 91.895 147.135 ;
        RECT 92.345 143.175 92.575 146.930 ;
        RECT 92.250 138.175 92.670 143.175 ;
        RECT 92.345 131.930 92.575 138.175 ;
        RECT 93.050 131.740 94.075 147.135 ;
        RECT 94.535 146.870 94.765 146.930 ;
        RECT 94.420 143.870 94.880 146.870 ;
        RECT 94.535 131.930 94.765 143.870 ;
        RECT 95.250 131.740 96.275 147.135 ;
        RECT 96.725 136.990 96.955 146.930 ;
        RECT 96.630 131.990 97.050 136.990 ;
        RECT 98.175 132.980 98.945 145.500 ;
        RECT 96.725 131.930 96.955 131.990 ;
        RECT 88.255 131.725 89.755 131.740 ;
        RECT 90.445 131.725 91.945 131.740 ;
        RECT 92.635 131.725 94.135 131.740 ;
        RECT 94.825 131.725 96.325 131.740 ;
        RECT 88.245 131.495 90.105 131.725 ;
        RECT 90.435 131.495 92.295 131.725 ;
        RECT 92.625 131.495 94.485 131.725 ;
        RECT 94.815 131.495 96.675 131.725 ;
        RECT 88.255 131.480 89.755 131.495 ;
        RECT 90.445 131.480 91.945 131.495 ;
        RECT 92.635 131.480 94.135 131.495 ;
        RECT 94.825 131.480 96.325 131.495 ;
        RECT 86.275 131.235 87.160 131.295 ;
        RECT 45.365 130.015 105.460 130.515 ;
        RECT 44.795 129.090 85.820 129.590 ;
        RECT 85.330 128.970 85.820 129.090 ;
        RECT 85.330 128.470 97.400 128.970 ;
        RECT 51.830 127.350 63.790 127.580 ;
        RECT 64.120 127.350 76.080 127.580 ;
        RECT 88.595 127.480 90.095 127.495 ;
        RECT 90.785 127.480 92.285 127.495 ;
        RECT 92.975 127.480 94.475 127.495 ;
        RECT 95.165 127.480 96.665 127.495 ;
        RECT 51.550 127.130 51.780 127.190 ;
        RECT 51.310 121.460 51.840 127.130 ;
        RECT 51.550 121.190 51.780 121.460 ;
        RECT 55.070 121.060 60.495 127.350 ;
        RECT 63.840 123.005 64.070 127.190 ;
        RECT 63.780 121.410 64.140 123.005 ;
        RECT 63.840 121.190 64.070 121.410 ;
        RECT 67.590 121.060 73.025 127.350 ;
        RECT 86.360 127.205 87.160 127.265 ;
        RECT 88.245 127.250 90.105 127.480 ;
        RECT 90.435 127.250 92.295 127.480 ;
        RECT 92.625 127.250 94.485 127.480 ;
        RECT 94.815 127.250 96.675 127.480 ;
        RECT 88.595 127.235 90.095 127.250 ;
        RECT 90.785 127.235 92.285 127.250 ;
        RECT 92.975 127.235 94.475 127.250 ;
        RECT 95.165 127.235 96.665 127.250 ;
        RECT 76.130 127.130 76.360 127.190 ;
        RECT 76.070 121.525 76.600 127.130 ;
        RECT 76.130 121.190 76.360 121.525 ;
        RECT 51.860 121.030 63.780 121.060 ;
        RECT 64.130 121.030 76.070 121.060 ;
        RECT 51.830 120.800 63.790 121.030 ;
        RECT 64.120 120.800 76.080 121.030 ;
        RECT 51.860 120.775 63.780 120.800 ;
        RECT 64.130 120.775 76.070 120.800 ;
        RECT 51.910 120.095 65.225 120.490 ;
        RECT 44.895 119.595 47.875 119.650 ;
        RECT 44.885 119.365 47.885 119.595 ;
        RECT 44.495 118.320 44.725 119.315 ;
        RECT 48.045 118.410 48.340 119.315 ;
        RECT 62.675 118.560 76.020 119.005 ;
        RECT 47.985 118.320 48.345 118.410 ;
        RECT 44.495 115.335 48.345 118.320 ;
        RECT 51.835 118.205 63.775 118.235 ;
        RECT 64.125 118.205 76.065 118.230 ;
        RECT 51.825 117.975 63.785 118.205 ;
        RECT 64.115 117.975 76.075 118.205 ;
        RECT 51.835 117.950 63.775 117.975 ;
        RECT 51.545 117.755 51.775 117.815 ;
        RECT 44.495 114.355 44.725 115.335 ;
        RECT 47.985 114.415 48.345 115.335 ;
        RECT 48.045 114.355 48.340 114.415 ;
        RECT 44.885 114.075 47.885 114.305 ;
        RECT 50.780 112.050 51.835 117.755 ;
        RECT 51.545 111.815 51.775 112.050 ;
        RECT 55.045 111.660 60.480 117.950 ;
        RECT 64.125 117.945 76.065 117.975 ;
        RECT 63.835 117.600 64.065 117.815 ;
        RECT 63.775 116.005 64.135 117.600 ;
        RECT 63.835 111.815 64.065 116.005 ;
        RECT 43.755 111.055 46.640 111.585 ;
        RECT 51.825 111.400 63.785 111.660 ;
        RECT 64.125 111.655 66.625 111.665 ;
        RECT 67.545 111.655 72.980 117.945 ;
        RECT 76.125 117.755 76.355 117.815 ;
        RECT 76.060 112.395 76.920 117.755 ;
        RECT 76.125 111.815 76.355 112.395 ;
        RECT 64.115 111.425 76.075 111.655 ;
        RECT 64.125 111.405 66.625 111.425 ;
        RECT 86.340 111.325 87.180 127.205 ;
        RECT 87.965 126.985 88.195 127.045 ;
        RECT 87.870 121.985 88.290 126.985 ;
        RECT 87.965 112.045 88.195 121.985 ;
        RECT 88.625 111.840 89.650 127.235 ;
        RECT 90.155 115.105 90.385 127.045 ;
        RECT 90.040 112.105 90.500 115.105 ;
        RECT 90.155 112.045 90.385 112.105 ;
        RECT 90.890 111.840 91.915 127.235 ;
        RECT 92.345 121.185 92.575 127.045 ;
        RECT 92.250 116.185 92.670 121.185 ;
        RECT 92.345 112.045 92.575 116.185 ;
        RECT 93.070 111.840 94.095 127.235 ;
        RECT 94.535 115.105 94.765 127.045 ;
        RECT 94.415 112.105 94.875 115.105 ;
        RECT 94.535 112.045 94.765 112.105 ;
        RECT 95.230 111.840 96.255 127.235 ;
        RECT 96.725 126.985 96.955 127.045 ;
        RECT 96.630 121.985 97.050 126.985 ;
        RECT 96.725 112.045 96.955 121.985 ;
        RECT 98.255 121.815 99.025 124.335 ;
        RECT 121.530 121.815 123.025 121.840 ;
        RECT 98.255 121.780 123.025 121.815 ;
        RECT 98.255 120.295 123.045 121.780 ;
        RECT 88.245 111.610 90.105 111.840 ;
        RECT 90.435 111.610 92.295 111.840 ;
        RECT 92.625 111.610 94.485 111.840 ;
        RECT 94.815 111.610 96.675 111.840 ;
        RECT 98.255 111.815 99.025 120.295 ;
        RECT 86.335 111.190 87.180 111.325 ;
        RECT 110.275 111.575 111.500 120.295 ;
        RECT 112.390 119.480 114.150 119.710 ;
        RECT 114.480 119.480 116.240 119.710 ;
        RECT 116.570 119.480 118.330 119.710 ;
        RECT 118.660 119.480 120.420 119.710 ;
        RECT 112.110 119.215 112.340 119.275 ;
        RECT 112.045 114.215 112.405 119.215 ;
        RECT 112.110 112.275 112.340 114.215 ;
        RECT 112.730 112.070 113.735 119.480 ;
        RECT 114.200 117.335 114.430 119.275 ;
        RECT 114.135 112.335 114.495 117.335 ;
        RECT 114.200 112.275 114.430 112.335 ;
        RECT 114.825 112.070 115.830 119.480 ;
        RECT 116.290 119.215 116.520 119.275 ;
        RECT 116.225 114.215 116.585 119.215 ;
        RECT 116.290 112.275 116.520 114.215 ;
        RECT 116.940 112.070 117.945 119.480 ;
        RECT 118.380 117.335 118.610 119.275 ;
        RECT 118.315 112.335 118.675 117.335 ;
        RECT 118.380 112.275 118.610 112.335 ;
        RECT 118.970 112.070 119.975 119.480 ;
        RECT 120.470 119.215 120.700 119.275 ;
        RECT 120.405 114.215 120.765 119.215 ;
        RECT 120.470 112.275 120.700 114.215 ;
        RECT 121.510 112.745 123.045 120.295 ;
        RECT 125.850 119.960 126.340 120.020 ;
        RECT 125.830 114.215 126.360 119.960 ;
        RECT 127.665 119.940 128.120 120.000 ;
        RECT 126.850 119.120 127.100 119.180 ;
        RECT 126.765 118.520 127.185 119.120 ;
        RECT 126.850 117.075 127.100 118.520 ;
        RECT 126.850 114.740 127.100 116.185 ;
        RECT 125.850 114.155 126.340 114.215 ;
        RECT 126.760 114.140 127.180 114.740 ;
        RECT 126.850 114.080 127.100 114.140 ;
        RECT 121.530 112.685 123.025 112.745 ;
        RECT 121.445 112.070 122.165 112.115 ;
        RECT 112.390 111.840 122.165 112.070 ;
        RECT 121.445 111.820 122.165 111.840 ;
        RECT 86.335 110.445 99.270 111.190 ;
        RECT 86.355 110.410 99.270 110.445 ;
        RECT 43.765 109.905 78.555 110.410 ;
        RECT 86.355 110.385 87.160 110.410 ;
        RECT 110.275 110.335 121.105 111.575 ;
        RECT 110.275 110.315 111.500 110.335 ;
        RECT 86.635 108.750 87.430 108.810 ;
        RECT 86.615 108.740 87.450 108.750 ;
        RECT 86.615 108.735 88.105 108.740 ;
        RECT 125.765 108.735 126.405 113.795 ;
        RECT 127.645 113.395 128.140 119.940 ;
        RECT 127.665 113.335 128.120 113.395 ;
        RECT 86.615 108.160 126.405 108.735 ;
        RECT 86.615 102.270 87.450 108.160 ;
        RECT 125.765 108.070 126.405 108.160 ;
        RECT 88.295 107.075 97.655 107.305 ;
        RECT 97.985 107.075 117.035 107.305 ;
        RECT 117.365 107.075 126.725 107.305 ;
        RECT 88.015 106.855 88.245 106.915 ;
        RECT 87.920 106.355 88.340 106.855 ;
        RECT 88.015 105.415 88.245 106.355 ;
        RECT 89.395 105.255 96.490 107.075 ;
        RECT 97.705 106.855 97.935 106.915 ;
        RECT 97.640 106.355 98.000 106.855 ;
        RECT 97.705 105.415 97.935 106.355 ;
        RECT 99.565 105.255 106.660 107.075 ;
        RECT 107.395 105.975 107.625 107.075 ;
        RECT 107.300 105.475 107.720 105.975 ;
        RECT 107.395 105.415 107.625 105.475 ;
        RECT 108.710 105.255 115.805 107.075 ;
        RECT 117.085 106.855 117.315 106.915 ;
        RECT 117.020 106.355 117.380 106.855 ;
        RECT 117.085 105.415 117.315 106.355 ;
        RECT 118.560 105.255 125.655 107.075 ;
        RECT 126.775 106.855 127.005 106.915 ;
        RECT 126.680 106.355 127.100 106.855 ;
        RECT 126.775 105.415 127.005 106.355 ;
        RECT 88.295 105.025 126.725 105.255 ;
        RECT 88.015 103.925 88.245 104.865 ;
        RECT 87.920 103.425 88.340 103.925 ;
        RECT 88.015 103.205 88.245 103.425 ;
        RECT 89.415 103.205 96.510 105.025 ;
        RECT 97.705 103.925 97.935 104.865 ;
        RECT 97.640 103.425 98.000 103.925 ;
        RECT 97.705 103.365 97.935 103.425 ;
        RECT 99.545 103.205 106.640 105.025 ;
        RECT 107.395 104.805 107.625 104.865 ;
        RECT 107.300 104.305 107.720 104.805 ;
        RECT 107.395 103.365 107.625 104.305 ;
        RECT 108.710 103.205 115.805 105.025 ;
        RECT 117.085 103.925 117.315 104.865 ;
        RECT 117.020 103.425 117.380 103.925 ;
        RECT 117.085 103.365 117.315 103.425 ;
        RECT 118.560 103.205 125.655 105.025 ;
        RECT 126.775 103.925 127.005 104.865 ;
        RECT 126.680 103.425 127.100 103.925 ;
        RECT 126.775 103.205 127.005 103.425 ;
        RECT 88.015 102.975 97.655 103.205 ;
        RECT 97.985 102.975 107.345 103.205 ;
        RECT 107.675 102.975 117.035 103.205 ;
        RECT 117.365 102.975 127.005 103.205 ;
        RECT 86.605 102.265 87.930 102.270 ;
        RECT 86.605 101.220 126.320 102.265 ;
        RECT 86.675 98.240 86.965 98.260 ;
        RECT 80.280 97.485 105.425 98.240 ;
        RECT 107.610 97.980 117.625 98.780 ;
        RECT 107.615 97.645 112.665 97.650 ;
        RECT 86.675 97.465 86.965 97.485 ;
        RECT 107.615 96.925 117.630 97.645 ;
        RECT 107.615 96.915 112.665 96.925 ;
        RECT 80.865 96.425 82.825 96.655 ;
        RECT 83.770 96.425 85.730 96.655 ;
        RECT 90.220 96.425 92.180 96.655 ;
        RECT 96.670 96.425 98.630 96.655 ;
        RECT 103.120 96.425 105.080 96.655 ;
        RECT 108.560 96.425 109.520 96.655 ;
        RECT 109.850 96.425 110.810 96.655 ;
        RECT 80.585 95.895 80.815 96.220 ;
        RECT 80.520 95.280 80.880 95.895 ;
        RECT 80.585 95.220 80.815 95.280 ;
        RECT 81.110 95.015 82.505 96.425 ;
        RECT 82.875 96.160 83.105 96.220 ;
        RECT 82.810 95.545 83.170 96.160 ;
        RECT 83.490 95.895 83.720 96.220 ;
        RECT 82.875 95.220 83.105 95.545 ;
        RECT 83.425 95.280 83.785 95.895 ;
        RECT 83.490 95.220 83.720 95.280 ;
        RECT 83.990 95.015 85.385 96.425 ;
        RECT 85.780 96.160 86.010 96.220 ;
        RECT 85.715 95.540 86.075 96.160 ;
        RECT 89.940 95.845 90.170 96.220 ;
        RECT 85.780 95.220 86.010 95.540 ;
        RECT 89.875 95.280 90.235 95.845 ;
        RECT 89.940 95.220 90.170 95.280 ;
        RECT 90.540 95.015 91.935 96.425 ;
        RECT 92.230 96.160 92.460 96.220 ;
        RECT 92.165 95.545 92.525 96.160 ;
        RECT 96.390 95.845 96.620 96.220 ;
        RECT 92.230 95.220 92.460 95.545 ;
        RECT 96.325 95.280 96.685 95.845 ;
        RECT 96.390 95.220 96.620 95.280 ;
        RECT 96.945 95.015 98.340 96.425 ;
        RECT 98.680 96.160 98.910 96.220 ;
        RECT 98.615 95.545 98.975 96.160 ;
        RECT 102.840 95.845 103.070 96.220 ;
        RECT 98.680 95.220 98.910 95.545 ;
        RECT 102.775 95.280 103.135 95.845 ;
        RECT 102.840 95.220 103.070 95.280 ;
        RECT 103.435 95.015 104.830 96.425 ;
        RECT 105.130 96.160 105.360 96.220 ;
        RECT 105.065 95.545 105.425 96.160 ;
        RECT 108.280 95.980 108.510 96.220 ;
        RECT 105.130 95.220 105.360 95.545 ;
        RECT 108.185 95.280 108.605 95.980 ;
        RECT 108.280 95.220 108.510 95.280 ;
        RECT 108.745 95.015 109.335 96.425 ;
        RECT 109.570 96.160 109.800 96.220 ;
        RECT 109.505 95.460 109.865 96.160 ;
        RECT 109.570 95.220 109.800 95.460 ;
        RECT 110.005 95.015 110.595 96.425 ;
        RECT 110.860 95.980 111.090 96.220 ;
        RECT 110.765 95.280 111.185 95.980 ;
        RECT 112.185 95.925 114.145 96.155 ;
        RECT 114.475 95.925 116.435 96.155 ;
        RECT 110.860 95.220 111.090 95.280 ;
        RECT 111.905 95.015 112.135 95.720 ;
        RECT 112.495 95.015 113.905 95.925 ;
        RECT 114.195 95.660 114.425 95.720 ;
        RECT 114.130 95.280 114.490 95.660 ;
        RECT 114.195 95.220 114.425 95.280 ;
        RECT 114.730 95.015 116.140 95.925 ;
        RECT 116.485 95.015 116.715 95.720 ;
        RECT 80.840 94.785 116.715 95.015 ;
        RECT 112.225 94.680 114.120 94.785 ;
        RECT 114.495 94.680 116.390 94.785 ;
        RECT 111.205 92.750 111.805 92.810 ;
        RECT 81.190 92.445 87.310 92.675 ;
        RECT 87.640 92.445 93.760 92.675 ;
        RECT 94.090 92.445 100.210 92.675 ;
        RECT 100.540 92.445 106.660 92.675 ;
        RECT 80.910 92.225 81.140 92.285 ;
        RECT 80.845 91.925 81.205 92.225 ;
        RECT 80.910 91.645 81.140 91.925 ;
        RECT 80.845 91.345 81.205 91.645 ;
        RECT 80.910 91.285 81.140 91.345 ;
        RECT 81.460 91.125 81.795 92.445 ;
        RECT 82.135 91.925 82.495 92.445 ;
        RECT 82.200 91.125 82.430 91.925 ;
        RECT 82.795 91.125 83.130 92.445 ;
        RECT 83.490 91.645 83.720 92.285 ;
        RECT 83.425 91.345 83.785 91.645 ;
        RECT 83.490 91.285 83.720 91.345 ;
        RECT 84.090 91.125 84.425 92.445 ;
        RECT 84.715 91.925 85.075 92.445 ;
        RECT 84.780 91.125 85.010 91.925 ;
        RECT 85.390 91.125 85.725 92.445 ;
        RECT 86.070 91.645 86.300 92.285 ;
        RECT 86.005 91.345 86.365 91.645 ;
        RECT 86.070 91.285 86.300 91.345 ;
        RECT 86.700 91.125 87.035 92.445 ;
        RECT 87.360 91.645 87.590 92.285 ;
        RECT 87.295 91.345 87.655 91.645 ;
        RECT 87.360 91.285 87.590 91.345 ;
        RECT 88.000 91.125 88.335 92.445 ;
        RECT 88.585 91.925 88.945 92.445 ;
        RECT 88.650 91.125 88.880 91.925 ;
        RECT 89.250 91.125 89.585 92.445 ;
        RECT 89.940 91.645 90.170 92.285 ;
        RECT 89.875 91.345 90.235 91.645 ;
        RECT 89.940 91.285 90.170 91.345 ;
        RECT 90.545 91.125 90.880 92.445 ;
        RECT 91.165 91.925 91.525 92.445 ;
        RECT 91.230 91.125 91.460 91.925 ;
        RECT 91.850 91.125 92.185 92.445 ;
        RECT 92.520 91.645 92.750 92.285 ;
        RECT 92.455 91.345 92.815 91.645 ;
        RECT 92.520 91.285 92.750 91.345 ;
        RECT 93.135 91.125 93.470 92.445 ;
        RECT 93.810 91.645 94.040 92.285 ;
        RECT 93.745 91.345 94.105 91.645 ;
        RECT 93.810 91.285 94.040 91.345 ;
        RECT 94.425 91.125 94.760 92.445 ;
        RECT 95.035 91.925 95.395 92.445 ;
        RECT 95.100 91.125 95.330 91.925 ;
        RECT 95.735 91.125 96.070 92.445 ;
        RECT 96.390 91.645 96.620 92.285 ;
        RECT 96.325 91.345 96.685 91.645 ;
        RECT 96.390 91.285 96.620 91.345 ;
        RECT 97.000 91.125 97.335 92.445 ;
        RECT 97.615 91.925 97.975 92.445 ;
        RECT 97.680 91.125 97.910 91.925 ;
        RECT 98.305 91.125 98.640 92.445 ;
        RECT 98.970 91.645 99.200 92.285 ;
        RECT 98.905 91.345 99.265 91.645 ;
        RECT 98.970 91.285 99.200 91.345 ;
        RECT 99.575 91.125 99.910 92.445 ;
        RECT 100.260 91.645 100.490 92.285 ;
        RECT 100.195 91.345 100.555 91.645 ;
        RECT 100.260 91.285 100.490 91.345 ;
        RECT 100.835 91.125 101.170 92.445 ;
        RECT 101.485 91.925 101.845 92.445 ;
        RECT 101.550 91.125 101.780 91.925 ;
        RECT 102.135 91.125 102.470 92.445 ;
        RECT 102.840 91.645 103.070 92.285 ;
        RECT 102.775 91.345 103.135 91.645 ;
        RECT 102.840 91.285 103.070 91.345 ;
        RECT 103.420 91.125 103.755 92.445 ;
        RECT 104.065 91.925 104.425 92.445 ;
        RECT 104.130 91.125 104.360 91.925 ;
        RECT 104.730 91.125 105.065 92.445 ;
        RECT 105.420 91.645 105.650 92.285 ;
        RECT 105.355 91.345 105.715 91.645 ;
        RECT 105.420 91.285 105.650 91.345 ;
        RECT 106.020 91.125 106.355 92.445 ;
        RECT 106.710 91.645 106.940 92.285 ;
        RECT 106.645 91.345 107.005 91.645 ;
        RECT 106.710 91.285 106.940 91.345 ;
        RECT 81.190 90.895 87.310 91.125 ;
        RECT 87.640 90.895 93.760 91.125 ;
        RECT 94.090 90.895 100.210 91.125 ;
        RECT 100.540 90.895 106.660 91.125 ;
        RECT 80.420 89.515 107.575 90.530 ;
        RECT 111.185 87.535 111.825 92.750 ;
        RECT 112.340 92.555 116.585 93.355 ;
        RECT 116.380 92.095 117.040 92.155 ;
        RECT 112.550 89.000 115.600 91.790 ;
        RECT 116.360 89.700 117.060 92.095 ;
        RECT 116.380 89.640 117.040 89.700 ;
        RECT 112.550 88.740 116.770 89.000 ;
        RECT 111.205 87.475 111.805 87.535 ;
        RECT 113.585 86.610 116.340 87.150 ;
        RECT 84.475 85.805 116.305 86.425 ;
        RECT 85.215 84.760 86.175 84.990 ;
        RECT 86.505 84.760 91.335 84.990 ;
        RECT 91.665 84.760 93.915 84.990 ;
        RECT 94.245 84.760 99.075 84.990 ;
        RECT 99.405 84.760 101.655 84.990 ;
        RECT 101.985 84.760 106.815 84.990 ;
        RECT 107.145 84.760 109.395 84.990 ;
        RECT 109.725 84.760 114.555 84.990 ;
        RECT 114.885 84.760 115.845 84.990 ;
        RECT 84.935 84.540 85.165 84.600 ;
        RECT 84.870 83.540 85.230 84.540 ;
        RECT 84.935 80.600 85.165 83.540 ;
        RECT 85.480 80.455 85.920 84.760 ;
        RECT 86.225 82.665 86.455 84.600 ;
        RECT 86.160 82.165 86.520 82.665 ;
        RECT 86.225 80.600 86.455 82.165 ;
        RECT 86.745 80.455 87.185 84.760 ;
        RECT 87.515 84.540 87.745 84.600 ;
        RECT 87.440 83.540 87.820 84.540 ;
        RECT 87.515 80.600 87.745 83.540 ;
        RECT 85.225 80.440 85.920 80.455 ;
        RECT 86.515 80.440 87.535 80.455 ;
        RECT 88.045 80.440 88.485 84.760 ;
        RECT 88.805 81.660 89.035 84.600 ;
        RECT 88.710 80.660 89.130 81.660 ;
        RECT 88.805 80.600 89.035 80.660 ;
        RECT 89.340 80.440 89.780 84.760 ;
        RECT 90.095 84.540 90.325 84.600 ;
        RECT 90.020 83.540 90.400 84.540 ;
        RECT 90.095 80.600 90.325 83.540 ;
        RECT 90.620 80.440 91.060 84.760 ;
        RECT 91.385 82.665 91.615 84.600 ;
        RECT 91.320 82.165 91.680 82.665 ;
        RECT 91.385 80.600 91.615 82.165 ;
        RECT 91.880 80.455 92.410 84.760 ;
        RECT 92.675 84.540 92.905 84.600 ;
        RECT 92.610 83.540 92.970 84.540 ;
        RECT 92.675 80.600 92.905 83.540 ;
        RECT 91.675 80.440 92.410 80.455 ;
        RECT 93.155 80.440 93.685 84.760 ;
        RECT 93.965 82.665 94.195 84.600 ;
        RECT 93.900 82.165 94.260 82.665 ;
        RECT 93.965 80.600 94.195 82.165 ;
        RECT 94.520 80.455 94.960 84.760 ;
        RECT 95.255 84.540 95.485 84.600 ;
        RECT 95.180 83.540 95.560 84.540 ;
        RECT 95.255 80.600 95.485 83.540 ;
        RECT 94.255 80.440 95.275 80.455 ;
        RECT 95.795 80.440 96.235 84.760 ;
        RECT 96.545 81.660 96.775 84.600 ;
        RECT 96.450 80.660 96.870 81.660 ;
        RECT 96.545 80.600 96.775 80.660 ;
        RECT 97.100 80.440 97.540 84.760 ;
        RECT 97.835 84.540 98.065 84.600 ;
        RECT 97.760 83.540 98.140 84.540 ;
        RECT 97.835 80.600 98.065 83.540 ;
        RECT 98.380 80.440 98.820 84.760 ;
        RECT 99.125 82.660 99.355 84.600 ;
        RECT 99.060 82.160 99.420 82.660 ;
        RECT 99.125 80.600 99.355 82.160 ;
        RECT 99.725 80.455 100.130 84.760 ;
        RECT 100.415 84.540 100.645 84.600 ;
        RECT 100.350 83.540 100.710 84.540 ;
        RECT 100.415 80.600 100.645 83.540 ;
        RECT 99.415 80.440 100.130 80.455 ;
        RECT 101.025 80.440 101.430 84.760 ;
        RECT 101.705 82.665 101.935 84.600 ;
        RECT 101.640 82.165 102.000 82.665 ;
        RECT 101.705 80.600 101.935 82.165 ;
        RECT 102.220 80.455 102.660 84.760 ;
        RECT 102.995 84.540 103.225 84.600 ;
        RECT 102.920 83.540 103.300 84.540 ;
        RECT 102.995 80.600 103.225 83.540 ;
        RECT 101.995 80.440 103.015 80.455 ;
        RECT 103.575 80.440 104.015 84.760 ;
        RECT 104.285 81.660 104.515 84.600 ;
        RECT 104.190 80.660 104.610 81.660 ;
        RECT 104.285 80.600 104.515 80.660 ;
        RECT 104.835 80.440 105.275 84.760 ;
        RECT 105.575 84.540 105.805 84.600 ;
        RECT 105.500 83.540 105.880 84.540 ;
        RECT 105.575 80.600 105.805 83.540 ;
        RECT 106.100 80.440 106.540 84.760 ;
        RECT 106.865 82.665 107.095 84.600 ;
        RECT 106.800 82.165 107.160 82.665 ;
        RECT 106.865 80.600 107.095 82.165 ;
        RECT 107.435 80.455 107.875 84.760 ;
        RECT 108.155 84.540 108.385 84.600 ;
        RECT 108.090 83.540 108.450 84.540 ;
        RECT 108.155 80.600 108.385 83.540 ;
        RECT 107.155 80.440 107.875 80.455 ;
        RECT 108.705 80.440 109.145 84.760 ;
        RECT 109.445 82.665 109.675 84.600 ;
        RECT 109.380 82.165 109.740 82.665 ;
        RECT 109.445 80.600 109.675 82.165 ;
        RECT 110.020 80.455 110.460 84.760 ;
        RECT 110.735 84.540 110.965 84.600 ;
        RECT 110.660 83.540 111.040 84.540 ;
        RECT 110.735 80.600 110.965 83.540 ;
        RECT 109.735 80.440 110.835 80.455 ;
        RECT 111.265 80.440 111.705 84.760 ;
        RECT 112.025 81.660 112.255 84.600 ;
        RECT 111.930 80.660 112.350 81.660 ;
        RECT 112.025 80.600 112.255 80.660 ;
        RECT 112.615 80.440 113.055 84.760 ;
        RECT 113.315 84.535 113.545 84.600 ;
        RECT 113.240 83.535 113.620 84.535 ;
        RECT 113.315 80.600 113.545 83.535 ;
        RECT 113.860 80.440 114.300 84.760 ;
        RECT 114.605 82.665 114.835 84.600 ;
        RECT 114.540 82.165 114.900 82.665 ;
        RECT 114.605 80.600 114.835 82.165 ;
        RECT 115.120 80.455 115.560 84.760 ;
        RECT 115.895 84.540 116.125 84.600 ;
        RECT 115.830 83.540 116.190 84.540 ;
        RECT 115.895 80.600 116.125 83.540 ;
        RECT 114.895 80.440 115.560 80.455 ;
        RECT 85.215 80.210 86.175 80.440 ;
        RECT 86.505 80.210 91.335 80.440 ;
        RECT 91.665 80.210 93.915 80.440 ;
        RECT 94.245 80.210 99.075 80.440 ;
        RECT 99.405 80.210 101.655 80.440 ;
        RECT 101.985 80.210 106.815 80.440 ;
        RECT 107.145 80.210 109.395 80.440 ;
        RECT 109.725 80.210 114.555 80.440 ;
        RECT 114.885 80.210 115.845 80.440 ;
        RECT 85.225 80.195 85.825 80.210 ;
        RECT 86.515 80.195 87.535 80.210 ;
        RECT 91.675 80.195 92.275 80.210 ;
        RECT 94.255 80.195 95.275 80.210 ;
        RECT 99.415 80.195 100.015 80.210 ;
        RECT 101.995 80.195 103.015 80.210 ;
        RECT 107.155 80.195 107.755 80.210 ;
        RECT 109.735 80.195 110.835 80.210 ;
        RECT 114.895 80.195 115.495 80.210 ;
        RECT 84.985 79.195 115.815 79.455 ;
        RECT 116.510 78.730 116.770 88.740 ;
        RECT 84.985 78.470 116.770 78.730 ;
        RECT 116.890 78.100 117.220 78.160 ;
        RECT 106.435 77.600 106.660 77.650 ;
        RECT 85.225 77.585 85.825 77.600 ;
        RECT 87.805 77.585 88.405 77.600 ;
        RECT 90.385 77.585 91.090 77.600 ;
        RECT 95.545 77.585 96.145 77.600 ;
        RECT 98.125 77.585 98.875 77.600 ;
        RECT 103.285 77.585 103.885 77.600 ;
        RECT 105.865 77.585 106.660 77.600 ;
        RECT 111.025 77.585 111.625 77.600 ;
        RECT 113.605 77.585 114.205 77.600 ;
        RECT 85.215 77.355 87.465 77.585 ;
        RECT 87.795 77.355 90.045 77.585 ;
        RECT 90.375 77.355 95.205 77.585 ;
        RECT 95.535 77.355 97.785 77.585 ;
        RECT 98.115 77.355 102.945 77.585 ;
        RECT 103.275 77.355 105.525 77.585 ;
        RECT 105.855 77.355 110.685 77.585 ;
        RECT 111.015 77.355 113.265 77.585 ;
        RECT 113.595 77.355 115.845 77.585 ;
        RECT 116.870 77.360 117.240 78.100 ;
        RECT 85.225 77.340 85.910 77.355 ;
        RECT 84.935 74.255 85.165 77.195 ;
        RECT 84.840 73.255 85.260 74.255 ;
        RECT 84.935 73.195 85.165 73.255 ;
        RECT 85.470 73.035 85.910 77.340 ;
        RECT 86.225 77.135 86.455 77.195 ;
        RECT 86.150 76.135 86.530 77.135 ;
        RECT 86.225 73.195 86.455 76.135 ;
        RECT 86.685 73.035 87.125 77.355 ;
        RECT 87.805 77.340 88.495 77.355 ;
        RECT 87.515 75.515 87.745 77.195 ;
        RECT 87.450 75.015 87.810 75.515 ;
        RECT 87.515 73.195 87.745 75.015 ;
        RECT 88.055 73.035 88.495 77.340 ;
        RECT 88.805 74.255 89.035 77.195 ;
        RECT 88.740 73.255 89.100 74.255 ;
        RECT 88.805 73.195 89.035 73.255 ;
        RECT 89.340 73.035 89.780 77.355 ;
        RECT 90.385 77.340 91.110 77.355 ;
        RECT 90.095 75.515 90.325 77.195 ;
        RECT 90.030 75.015 90.390 75.515 ;
        RECT 90.095 73.195 90.325 75.015 ;
        RECT 90.670 73.035 91.110 77.340 ;
        RECT 91.385 77.135 91.615 77.195 ;
        RECT 91.310 76.135 91.690 77.135 ;
        RECT 91.385 73.195 91.615 76.135 ;
        RECT 91.925 73.035 92.365 77.355 ;
        RECT 92.675 74.255 92.905 77.195 ;
        RECT 92.580 73.255 93.000 74.255 ;
        RECT 92.675 73.195 92.905 73.255 ;
        RECT 93.250 73.035 93.690 77.355 ;
        RECT 93.965 77.135 94.195 77.195 ;
        RECT 93.890 76.135 94.270 77.135 ;
        RECT 93.965 73.195 94.195 76.135 ;
        RECT 94.470 73.035 94.910 77.355 ;
        RECT 95.545 77.340 96.245 77.355 ;
        RECT 95.255 75.515 95.485 77.195 ;
        RECT 95.190 75.015 95.550 75.515 ;
        RECT 95.255 73.195 95.485 75.015 ;
        RECT 95.805 73.035 96.245 77.340 ;
        RECT 96.545 74.255 96.775 77.195 ;
        RECT 96.485 73.255 96.845 74.255 ;
        RECT 96.545 73.195 96.775 73.255 ;
        RECT 97.090 73.035 97.530 77.355 ;
        RECT 98.125 77.340 98.875 77.355 ;
        RECT 97.835 75.515 98.065 77.195 ;
        RECT 97.770 75.015 98.130 75.515 ;
        RECT 97.835 73.195 98.065 75.015 ;
        RECT 98.350 73.035 98.790 77.340 ;
        RECT 99.125 77.135 99.355 77.195 ;
        RECT 99.050 76.135 99.430 77.135 ;
        RECT 99.125 73.195 99.355 76.135 ;
        RECT 99.645 73.035 100.085 77.355 ;
        RECT 100.415 74.255 100.645 77.195 ;
        RECT 100.320 73.255 100.740 74.255 ;
        RECT 100.415 73.195 100.645 73.255 ;
        RECT 100.930 73.035 101.370 77.355 ;
        RECT 101.705 77.135 101.935 77.195 ;
        RECT 101.630 76.135 102.010 77.135 ;
        RECT 101.705 73.195 101.935 76.135 ;
        RECT 102.210 73.035 102.650 77.355 ;
        RECT 103.285 77.340 103.975 77.355 ;
        RECT 102.995 75.515 103.225 77.195 ;
        RECT 102.930 75.015 103.290 75.515 ;
        RECT 102.995 73.195 103.225 75.015 ;
        RECT 103.535 73.035 103.975 77.340 ;
        RECT 104.285 74.255 104.515 77.195 ;
        RECT 104.220 73.255 104.580 74.255 ;
        RECT 104.285 73.195 104.515 73.255 ;
        RECT 104.820 73.035 105.285 77.355 ;
        RECT 105.865 77.340 106.660 77.355 ;
        RECT 106.110 77.290 106.660 77.340 ;
        RECT 105.575 75.515 105.805 77.195 ;
        RECT 105.510 75.015 105.870 75.515 ;
        RECT 105.575 73.195 105.805 75.015 ;
        RECT 106.110 73.035 106.550 77.290 ;
        RECT 106.865 77.135 107.095 77.195 ;
        RECT 106.790 76.135 107.170 77.135 ;
        RECT 106.865 73.195 107.095 76.135 ;
        RECT 107.405 73.035 107.845 77.355 ;
        RECT 108.155 74.255 108.385 77.195 ;
        RECT 108.060 73.255 108.480 74.255 ;
        RECT 108.155 73.195 108.385 73.255 ;
        RECT 108.655 73.035 109.095 77.355 ;
        RECT 109.445 77.135 109.675 77.195 ;
        RECT 109.370 76.135 109.750 77.135 ;
        RECT 109.445 73.195 109.675 76.135 ;
        RECT 109.970 73.035 110.410 77.355 ;
        RECT 111.025 77.340 111.715 77.355 ;
        RECT 110.735 75.515 110.965 77.195 ;
        RECT 110.670 75.015 111.030 75.515 ;
        RECT 110.735 73.195 110.965 75.015 ;
        RECT 111.275 73.035 111.715 77.340 ;
        RECT 112.025 74.255 112.255 77.195 ;
        RECT 111.960 73.255 112.320 74.255 ;
        RECT 112.025 73.195 112.255 73.255 ;
        RECT 112.590 73.035 113.035 77.355 ;
        RECT 113.605 77.340 114.280 77.355 ;
        RECT 113.315 75.515 113.545 77.195 ;
        RECT 113.250 75.015 113.610 75.515 ;
        RECT 113.315 73.195 113.545 75.015 ;
        RECT 113.835 73.035 114.280 77.340 ;
        RECT 114.605 77.135 114.835 77.195 ;
        RECT 114.530 76.135 114.910 77.135 ;
        RECT 114.605 73.195 114.835 76.135 ;
        RECT 115.155 73.035 115.600 77.355 ;
        RECT 116.890 77.300 117.220 77.360 ;
        RECT 115.895 74.255 116.125 77.195 ;
        RECT 115.800 73.255 116.220 74.255 ;
        RECT 115.895 73.195 116.125 73.255 ;
        RECT 116.890 73.170 117.220 73.230 ;
        RECT 85.215 72.805 87.465 73.035 ;
        RECT 87.795 72.805 90.045 73.035 ;
        RECT 90.375 72.805 95.205 73.035 ;
        RECT 95.535 72.805 97.785 73.035 ;
        RECT 98.115 72.805 102.945 73.035 ;
        RECT 103.275 72.805 105.525 73.035 ;
        RECT 105.855 72.805 110.685 73.035 ;
        RECT 111.015 72.805 113.265 73.035 ;
        RECT 113.595 72.805 115.845 73.035 ;
        RECT 116.870 72.410 117.240 73.170 ;
        RECT 116.890 72.350 117.220 72.410 ;
        RECT 84.255 71.100 117.265 72.030 ;
        RECT 89.490 55.045 128.600 55.550 ;
        RECT 90.140 53.535 127.375 53.765 ;
        RECT 13.410 19.085 14.340 52.095 ;
        RECT 14.720 52.050 15.480 52.070 ;
        RECT 19.670 52.050 20.410 52.070 ;
        RECT 14.660 51.720 15.540 52.050 ;
        RECT 19.610 51.720 20.470 52.050 ;
        RECT 32.010 51.870 34.405 51.890 ;
        RECT 14.720 51.700 15.480 51.720 ;
        RECT 19.670 51.700 20.410 51.720 ;
        RECT 20.780 51.340 31.310 51.600 ;
        RECT 15.565 50.955 16.565 51.050 ;
        RECT 15.505 50.725 19.505 50.955 ;
        RECT 15.115 50.430 15.345 50.675 ;
        RECT 15.565 50.630 16.565 50.725 ;
        RECT 19.665 50.430 19.895 50.675 ;
        RECT 15.115 49.985 19.895 50.430 ;
        RECT 15.115 49.110 15.345 49.985 ;
        RECT 18.445 49.665 19.445 49.740 ;
        RECT 15.505 49.435 19.505 49.665 ;
        RECT 18.445 49.360 19.445 49.435 ;
        RECT 19.665 49.110 19.895 49.985 ;
        RECT 15.115 49.035 19.895 49.110 ;
        RECT 15.115 48.665 19.910 49.035 ;
        RECT 15.115 48.425 15.345 48.665 ;
        RECT 17.325 48.375 17.825 48.440 ;
        RECT 19.650 48.435 19.910 48.665 ;
        RECT 19.665 48.425 19.895 48.435 ;
        RECT 15.505 48.145 19.505 48.375 ;
        RECT 15.115 47.865 15.345 48.095 ;
        RECT 17.325 48.080 17.825 48.145 ;
        RECT 19.665 47.865 19.895 48.095 ;
        RECT 15.115 47.420 19.895 47.865 ;
        RECT 15.115 46.545 15.345 47.420 ;
        RECT 15.565 47.085 16.565 47.150 ;
        RECT 15.505 46.855 19.505 47.085 ;
        RECT 15.565 46.790 16.565 46.855 ;
        RECT 19.665 46.545 19.895 47.420 ;
        RECT 15.115 46.455 19.895 46.545 ;
        RECT 15.115 46.105 19.910 46.455 ;
        RECT 15.115 45.845 15.345 46.105 ;
        RECT 17.325 45.795 17.825 45.860 ;
        RECT 19.650 45.855 19.910 46.105 ;
        RECT 19.665 45.845 19.895 45.855 ;
        RECT 15.505 45.565 19.505 45.795 ;
        RECT 15.115 45.240 15.345 45.515 ;
        RECT 17.325 45.500 17.825 45.565 ;
        RECT 19.665 45.240 19.895 45.515 ;
        RECT 15.115 44.800 19.895 45.240 ;
        RECT 15.115 43.925 15.345 44.800 ;
        RECT 18.445 44.505 19.445 44.580 ;
        RECT 15.505 44.275 19.505 44.505 ;
        RECT 18.445 44.200 19.445 44.275 ;
        RECT 19.665 43.925 19.895 44.800 ;
        RECT 15.115 43.485 19.895 43.925 ;
        RECT 15.115 42.675 15.345 43.485 ;
        RECT 15.565 43.215 16.565 43.310 ;
        RECT 15.505 42.985 19.505 43.215 ;
        RECT 15.565 42.890 16.565 42.985 ;
        RECT 19.665 42.675 19.895 43.485 ;
        RECT 15.115 42.235 19.895 42.675 ;
        RECT 15.115 41.380 15.345 42.235 ;
        RECT 18.445 41.925 19.445 42.000 ;
        RECT 15.505 41.695 19.505 41.925 ;
        RECT 18.445 41.620 19.445 41.695 ;
        RECT 19.665 41.490 19.895 42.235 ;
        RECT 19.600 41.380 19.960 41.490 ;
        RECT 15.115 41.265 19.960 41.380 ;
        RECT 15.115 40.940 19.910 41.265 ;
        RECT 15.115 40.685 15.345 40.940 ;
        RECT 17.325 40.635 17.825 40.700 ;
        RECT 19.650 40.695 19.910 40.940 ;
        RECT 19.665 40.685 19.895 40.695 ;
        RECT 15.505 40.405 19.505 40.635 ;
        RECT 15.115 40.115 15.345 40.355 ;
        RECT 17.325 40.340 17.825 40.405 ;
        RECT 19.665 40.115 19.895 40.355 ;
        RECT 15.115 39.650 19.895 40.115 ;
        RECT 15.115 38.805 15.345 39.650 ;
        RECT 15.565 39.345 16.565 39.410 ;
        RECT 15.505 39.115 19.505 39.345 ;
        RECT 15.565 39.050 16.565 39.115 ;
        RECT 19.665 38.805 19.895 39.650 ;
        RECT 15.115 38.715 19.895 38.805 ;
        RECT 15.115 38.365 19.910 38.715 ;
        RECT 15.115 38.105 15.345 38.365 ;
        RECT 17.325 38.055 17.825 38.120 ;
        RECT 19.650 38.115 19.910 38.365 ;
        RECT 19.665 38.105 19.895 38.115 ;
        RECT 15.505 37.825 19.505 38.055 ;
        RECT 15.115 37.480 15.345 37.775 ;
        RECT 17.325 37.760 17.825 37.825 ;
        RECT 19.665 37.480 19.895 37.775 ;
        RECT 15.115 37.040 19.895 37.480 ;
        RECT 15.115 36.200 15.345 37.040 ;
        RECT 18.445 36.765 19.445 36.840 ;
        RECT 15.505 36.535 19.505 36.765 ;
        RECT 18.445 36.460 19.445 36.535 ;
        RECT 19.665 36.200 19.895 37.040 ;
        RECT 15.115 35.760 19.895 36.200 ;
        RECT 15.115 34.915 15.345 35.760 ;
        RECT 15.565 35.475 16.565 35.570 ;
        RECT 15.505 35.245 19.505 35.475 ;
        RECT 15.565 35.150 16.565 35.245 ;
        RECT 19.665 34.915 19.895 35.760 ;
        RECT 15.115 34.475 19.895 34.915 ;
        RECT 15.115 33.620 15.345 34.475 ;
        RECT 18.445 34.185 19.445 34.260 ;
        RECT 15.505 33.955 19.505 34.185 ;
        RECT 18.445 33.880 19.445 33.955 ;
        RECT 19.665 33.705 19.895 34.475 ;
        RECT 19.650 33.620 19.910 33.705 ;
        RECT 15.115 33.180 19.910 33.620 ;
        RECT 15.115 32.945 15.345 33.180 ;
        RECT 17.325 32.895 17.825 32.960 ;
        RECT 19.650 32.955 19.910 33.180 ;
        RECT 19.665 32.945 19.895 32.955 ;
        RECT 15.505 32.665 19.505 32.895 ;
        RECT 15.115 32.360 15.345 32.615 ;
        RECT 17.325 32.600 17.825 32.665 ;
        RECT 19.665 32.360 19.895 32.615 ;
        RECT 15.115 31.920 19.895 32.360 ;
        RECT 15.115 31.075 15.345 31.920 ;
        RECT 15.565 31.605 16.565 31.675 ;
        RECT 15.505 31.375 19.505 31.605 ;
        RECT 15.565 31.315 16.565 31.375 ;
        RECT 19.665 31.075 19.895 31.920 ;
        RECT 15.115 30.975 19.895 31.075 ;
        RECT 15.115 30.635 19.910 30.975 ;
        RECT 15.115 30.365 15.345 30.635 ;
        RECT 17.325 30.315 17.825 30.380 ;
        RECT 19.650 30.375 19.910 30.635 ;
        RECT 19.665 30.365 19.895 30.375 ;
        RECT 15.505 30.085 19.505 30.315 ;
        RECT 15.115 29.740 15.345 30.035 ;
        RECT 17.325 30.020 17.825 30.085 ;
        RECT 19.665 29.740 19.895 30.035 ;
        RECT 15.115 29.300 19.895 29.740 ;
        RECT 15.115 28.520 15.345 29.300 ;
        RECT 18.445 29.025 19.445 29.100 ;
        RECT 15.505 28.795 19.505 29.025 ;
        RECT 18.445 28.720 19.445 28.795 ;
        RECT 19.665 28.520 19.895 29.300 ;
        RECT 15.115 28.080 19.895 28.520 ;
        RECT 15.115 27.195 15.345 28.080 ;
        RECT 15.565 27.735 16.565 27.830 ;
        RECT 15.505 27.505 19.505 27.735 ;
        RECT 15.565 27.410 16.565 27.505 ;
        RECT 19.665 27.195 19.895 28.080 ;
        RECT 15.115 26.755 19.895 27.195 ;
        RECT 15.115 25.940 15.345 26.755 ;
        RECT 18.445 26.445 19.445 26.520 ;
        RECT 15.505 26.215 19.505 26.445 ;
        RECT 18.445 26.140 19.445 26.215 ;
        RECT 19.665 25.940 19.895 26.755 ;
        RECT 15.115 25.920 19.895 25.940 ;
        RECT 15.115 25.500 19.910 25.920 ;
        RECT 15.115 25.205 15.345 25.500 ;
        RECT 17.325 25.155 17.825 25.220 ;
        RECT 19.650 25.215 19.910 25.500 ;
        RECT 19.665 25.205 19.895 25.215 ;
        RECT 15.505 24.925 19.505 25.155 ;
        RECT 15.115 24.610 15.345 24.875 ;
        RECT 17.325 24.860 17.825 24.925 ;
        RECT 19.665 24.610 19.895 24.875 ;
        RECT 15.115 24.170 19.895 24.610 ;
        RECT 15.115 23.325 15.345 24.170 ;
        RECT 15.565 23.865 16.565 23.930 ;
        RECT 15.505 23.635 19.505 23.865 ;
        RECT 15.565 23.570 16.565 23.635 ;
        RECT 19.665 23.325 19.895 24.170 ;
        RECT 15.115 23.235 19.895 23.325 ;
        RECT 15.115 22.885 19.910 23.235 ;
        RECT 15.115 22.625 15.345 22.885 ;
        RECT 17.325 22.575 17.825 22.640 ;
        RECT 19.650 22.635 19.910 22.885 ;
        RECT 19.665 22.625 19.895 22.635 ;
        RECT 15.505 22.345 19.505 22.575 ;
        RECT 15.115 21.955 15.345 22.295 ;
        RECT 17.325 22.280 17.825 22.345 ;
        RECT 19.665 21.955 19.895 22.295 ;
        RECT 15.115 21.515 19.895 21.955 ;
        RECT 15.115 20.740 15.345 21.515 ;
        RECT 18.445 21.285 19.445 21.360 ;
        RECT 15.505 21.055 19.505 21.285 ;
        RECT 18.445 20.980 19.445 21.055 ;
        RECT 19.665 20.740 19.895 21.515 ;
        RECT 15.115 20.655 19.895 20.740 ;
        RECT 15.115 20.300 19.910 20.655 ;
        RECT 15.115 20.045 15.345 20.300 ;
        RECT 15.565 19.995 16.565 20.090 ;
        RECT 19.650 20.055 19.910 20.300 ;
        RECT 19.665 20.045 19.895 20.055 ;
        RECT 15.505 19.765 19.505 19.995 ;
        RECT 20.780 19.815 21.040 51.340 ;
        RECT 25.850 50.955 26.850 51.020 ;
        RECT 22.910 50.725 26.910 50.955 ;
        RECT 21.505 19.815 21.765 50.645 ;
        RECT 22.520 50.390 22.750 50.675 ;
        RECT 25.850 50.660 26.850 50.725 ;
        RECT 27.070 50.390 27.300 50.675 ;
        RECT 22.520 50.325 27.300 50.390 ;
        RECT 22.505 49.950 27.300 50.325 ;
        RECT 22.505 49.725 22.765 49.950 ;
        RECT 22.520 49.715 22.750 49.725 ;
        RECT 24.475 49.665 24.975 49.730 ;
        RECT 27.070 49.715 27.300 49.950 ;
        RECT 22.910 49.435 26.910 49.665 ;
        RECT 22.520 49.130 22.750 49.385 ;
        RECT 24.475 49.370 24.975 49.435 ;
        RECT 27.070 49.130 27.300 49.385 ;
        RECT 22.520 48.690 27.300 49.130 ;
        RECT 22.520 47.885 22.750 48.690 ;
        RECT 25.845 48.375 26.845 48.450 ;
        RECT 22.910 48.145 26.910 48.375 ;
        RECT 25.845 48.070 26.845 48.145 ;
        RECT 27.070 47.885 27.300 48.690 ;
        RECT 22.520 47.445 27.300 47.885 ;
        RECT 22.520 46.535 22.750 47.445 ;
        RECT 22.970 47.085 23.970 47.180 ;
        RECT 22.910 46.855 26.910 47.085 ;
        RECT 22.970 46.760 23.970 46.855 ;
        RECT 27.070 46.535 27.300 47.445 ;
        RECT 22.520 46.095 27.300 46.535 ;
        RECT 22.520 45.665 22.750 46.095 ;
        RECT 25.850 45.795 26.850 45.870 ;
        RECT 22.505 45.290 22.765 45.665 ;
        RECT 22.910 45.565 26.910 45.795 ;
        RECT 25.850 45.490 26.850 45.565 ;
        RECT 27.070 45.290 27.300 46.095 ;
        RECT 22.505 44.850 27.300 45.290 ;
        RECT 22.505 44.565 22.765 44.850 ;
        RECT 22.520 44.555 22.750 44.565 ;
        RECT 24.475 44.505 24.975 44.570 ;
        RECT 27.070 44.555 27.300 44.850 ;
        RECT 22.910 44.275 26.910 44.505 ;
        RECT 22.520 43.975 22.750 44.225 ;
        RECT 24.475 44.210 24.975 44.275 ;
        RECT 27.070 43.975 27.300 44.225 ;
        RECT 22.520 43.535 27.300 43.975 ;
        RECT 22.520 42.705 22.750 43.535 ;
        RECT 25.850 43.215 26.850 43.280 ;
        RECT 22.910 42.985 26.910 43.215 ;
        RECT 25.850 42.920 26.850 42.985 ;
        RECT 27.070 42.705 27.300 43.535 ;
        RECT 22.520 42.585 27.300 42.705 ;
        RECT 22.505 42.265 27.300 42.585 ;
        RECT 22.505 41.985 22.765 42.265 ;
        RECT 22.520 41.975 22.750 41.985 ;
        RECT 24.475 41.925 24.975 41.990 ;
        RECT 27.070 41.975 27.300 42.265 ;
        RECT 22.910 41.695 26.910 41.925 ;
        RECT 22.520 41.370 22.750 41.645 ;
        RECT 24.475 41.630 24.975 41.695 ;
        RECT 27.070 41.370 27.300 41.645 ;
        RECT 22.520 40.930 27.300 41.370 ;
        RECT 22.520 40.105 22.750 40.930 ;
        RECT 25.850 40.635 26.850 40.710 ;
        RECT 22.910 40.405 26.910 40.635 ;
        RECT 25.850 40.330 26.850 40.405 ;
        RECT 27.070 40.105 27.300 40.930 ;
        RECT 22.520 39.665 27.300 40.105 ;
        RECT 22.520 38.845 22.750 39.665 ;
        RECT 22.970 39.345 23.970 39.440 ;
        RECT 22.910 39.115 26.910 39.345 ;
        RECT 22.970 39.020 23.970 39.115 ;
        RECT 27.070 38.845 27.300 39.665 ;
        RECT 22.520 38.405 27.300 38.845 ;
        RECT 22.520 37.845 22.750 38.405 ;
        RECT 25.850 38.055 26.850 38.130 ;
        RECT 22.505 37.490 22.765 37.845 ;
        RECT 22.910 37.825 26.910 38.055 ;
        RECT 25.850 37.750 26.850 37.825 ;
        RECT 27.070 37.490 27.300 38.405 ;
        RECT 22.505 37.050 27.300 37.490 ;
        RECT 22.505 36.825 22.765 37.050 ;
        RECT 22.520 36.815 22.750 36.825 ;
        RECT 24.475 36.765 24.975 36.830 ;
        RECT 27.070 36.815 27.300 37.050 ;
        RECT 22.910 36.535 26.910 36.765 ;
        RECT 22.520 36.260 22.750 36.485 ;
        RECT 24.475 36.470 24.975 36.535 ;
        RECT 27.070 36.260 27.300 36.485 ;
        RECT 22.520 35.855 27.300 36.260 ;
        RECT 22.520 34.960 22.750 35.855 ;
        RECT 25.850 35.475 26.850 35.540 ;
        RECT 22.910 35.245 26.910 35.475 ;
        RECT 25.850 35.180 26.850 35.245 ;
        RECT 27.070 34.960 27.300 35.855 ;
        RECT 22.520 34.845 27.300 34.960 ;
        RECT 22.505 34.555 27.300 34.845 ;
        RECT 22.505 34.245 22.765 34.555 ;
        RECT 22.520 34.235 22.750 34.245 ;
        RECT 24.470 34.185 24.970 34.250 ;
        RECT 27.070 34.235 27.300 34.555 ;
        RECT 22.910 33.955 26.910 34.185 ;
        RECT 22.520 33.650 22.750 33.905 ;
        RECT 24.470 33.890 24.970 33.955 ;
        RECT 27.070 33.650 27.300 33.905 ;
        RECT 22.520 33.210 27.300 33.650 ;
        RECT 22.520 32.370 22.750 33.210 ;
        RECT 25.850 32.895 26.850 32.970 ;
        RECT 22.910 32.665 26.910 32.895 ;
        RECT 25.850 32.590 26.850 32.665 ;
        RECT 27.070 32.370 27.300 33.210 ;
        RECT 22.520 31.930 27.300 32.370 ;
        RECT 22.520 31.065 22.750 31.930 ;
        RECT 22.970 31.605 23.970 31.700 ;
        RECT 22.910 31.375 26.910 31.605 ;
        RECT 22.970 31.280 23.970 31.375 ;
        RECT 27.070 31.065 27.300 31.930 ;
        RECT 22.520 30.625 27.300 31.065 ;
        RECT 22.520 30.105 22.750 30.625 ;
        RECT 25.850 30.315 26.850 30.390 ;
        RECT 22.505 29.790 22.765 30.105 ;
        RECT 22.910 30.085 26.910 30.315 ;
        RECT 25.850 30.010 26.850 30.085 ;
        RECT 27.070 29.790 27.300 30.625 ;
        RECT 22.505 29.350 27.300 29.790 ;
        RECT 22.505 29.085 22.765 29.350 ;
        RECT 22.520 29.075 22.750 29.085 ;
        RECT 24.475 29.025 24.975 29.090 ;
        RECT 27.070 29.075 27.300 29.350 ;
        RECT 22.910 28.795 26.910 29.025 ;
        RECT 22.520 28.515 22.750 28.745 ;
        RECT 24.475 28.730 24.975 28.795 ;
        RECT 27.070 28.515 27.300 28.745 ;
        RECT 22.520 27.985 27.300 28.515 ;
        RECT 22.520 27.240 22.750 27.985 ;
        RECT 25.850 27.735 26.850 27.800 ;
        RECT 22.910 27.505 26.910 27.735 ;
        RECT 25.850 27.440 26.850 27.505 ;
        RECT 27.070 27.240 27.300 27.985 ;
        RECT 22.520 27.105 27.300 27.240 ;
        RECT 22.505 26.710 27.300 27.105 ;
        RECT 22.505 26.505 22.765 26.710 ;
        RECT 22.520 26.495 22.750 26.505 ;
        RECT 24.475 26.445 24.975 26.510 ;
        RECT 27.070 26.495 27.300 26.710 ;
        RECT 22.910 26.215 26.910 26.445 ;
        RECT 22.520 25.890 22.750 26.165 ;
        RECT 24.475 26.150 24.975 26.215 ;
        RECT 27.070 25.890 27.300 26.165 ;
        RECT 22.520 25.450 27.300 25.890 ;
        RECT 22.520 24.610 22.750 25.450 ;
        RECT 25.850 25.155 26.850 25.230 ;
        RECT 22.910 24.925 26.910 25.155 ;
        RECT 25.850 24.850 26.850 24.925 ;
        RECT 27.070 24.610 27.300 25.450 ;
        RECT 22.520 24.170 27.300 24.610 ;
        RECT 22.520 23.315 22.750 24.170 ;
        RECT 22.970 23.865 23.970 23.960 ;
        RECT 22.910 23.635 26.910 23.865 ;
        RECT 22.970 23.540 23.970 23.635 ;
        RECT 27.070 23.315 27.300 24.170 ;
        RECT 22.520 22.875 27.300 23.315 ;
        RECT 22.520 22.365 22.750 22.875 ;
        RECT 25.850 22.575 26.850 22.650 ;
        RECT 22.505 22.015 22.765 22.365 ;
        RECT 22.910 22.345 26.910 22.575 ;
        RECT 25.850 22.270 26.850 22.345 ;
        RECT 27.070 22.015 27.300 22.875 ;
        RECT 22.505 21.575 27.300 22.015 ;
        RECT 22.505 21.345 22.765 21.575 ;
        RECT 22.520 21.335 22.750 21.345 ;
        RECT 24.475 21.285 24.975 21.350 ;
        RECT 27.070 21.335 27.300 21.575 ;
        RECT 22.910 21.055 26.910 21.285 ;
        RECT 22.520 20.750 22.750 21.005 ;
        RECT 24.475 20.990 24.975 21.055 ;
        RECT 27.070 20.750 27.300 21.005 ;
        RECT 22.520 20.655 27.300 20.750 ;
        RECT 22.505 20.310 27.300 20.655 ;
        RECT 22.505 20.055 22.765 20.310 ;
        RECT 22.520 20.045 22.750 20.055 ;
        RECT 25.850 19.995 26.850 20.060 ;
        RECT 27.070 20.045 27.300 20.310 ;
        RECT 22.910 19.765 26.910 19.995 ;
        RECT 15.565 19.670 16.565 19.765 ;
        RECT 25.850 19.700 26.850 19.765 ;
        RECT 28.115 19.305 28.735 51.135 ;
        RECT 28.920 48.415 29.460 51.170 ;
        RECT 31.050 50.430 31.310 51.340 ;
        RECT 31.950 51.210 34.465 51.870 ;
        RECT 32.010 51.190 34.405 51.210 ;
        RECT 31.050 47.380 34.100 50.430 ;
        RECT 34.865 47.170 35.665 51.415 ;
        RECT 37.095 51.315 38.030 51.545 ;
        RECT 37.095 51.220 37.325 51.315 ;
        RECT 36.990 50.970 37.325 51.220 ;
        RECT 38.235 50.970 38.465 51.265 ;
        RECT 36.990 49.560 38.465 50.970 ;
        RECT 36.990 49.325 37.325 49.560 ;
        RECT 37.095 48.950 37.325 49.325 ;
        RECT 37.590 49.255 37.970 49.320 ;
        RECT 38.235 49.305 38.465 49.560 ;
        RECT 37.530 49.025 38.030 49.255 ;
        RECT 37.590 48.960 37.970 49.025 ;
        RECT 36.990 48.735 37.325 48.950 ;
        RECT 38.235 48.735 38.465 48.975 ;
        RECT 36.990 47.325 38.465 48.735 ;
        RECT 39.235 47.495 39.955 52.460 ;
        RECT 36.990 47.055 37.325 47.325 ;
        RECT 37.095 46.965 37.325 47.055 ;
        RECT 38.235 47.015 38.465 47.325 ;
        RECT 37.095 46.735 38.030 46.965 ;
        RECT 29.845 46.635 35.060 46.655 ;
        RECT 29.785 46.035 35.120 46.635 ;
        RECT 29.845 46.015 35.060 46.035 ;
        RECT 37.095 45.425 37.325 46.735 ;
        RECT 37.590 45.920 38.290 46.015 ;
        RECT 37.530 45.690 38.530 45.920 ;
        RECT 37.590 45.595 38.290 45.690 ;
        RECT 38.735 45.425 38.965 45.640 ;
        RECT 37.095 44.835 38.965 45.425 ;
        RECT 37.095 44.165 37.325 44.835 ;
        RECT 37.770 44.630 38.470 44.695 ;
        RECT 38.735 44.680 38.965 44.835 ;
        RECT 37.530 44.400 38.530 44.630 ;
        RECT 37.770 44.335 38.470 44.400 ;
        RECT 38.735 44.165 38.965 44.350 ;
        RECT 37.095 43.575 38.965 44.165 ;
        RECT 31.825 14.755 32.840 41.910 ;
        RECT 33.655 41.275 33.955 41.340 ;
        RECT 33.595 41.045 34.595 41.275 ;
        RECT 33.205 40.690 33.435 40.995 ;
        RECT 33.655 40.980 33.955 41.045 ;
        RECT 34.755 40.690 34.985 40.995 ;
        RECT 33.205 40.355 34.985 40.690 ;
        RECT 33.205 39.400 33.435 40.355 ;
        RECT 33.655 39.985 33.955 40.050 ;
        RECT 33.595 39.755 34.595 39.985 ;
        RECT 33.655 39.690 33.955 39.755 ;
        RECT 34.755 39.400 34.985 40.355 ;
        RECT 33.205 39.065 34.985 39.400 ;
        RECT 33.205 38.695 33.435 39.065 ;
        RECT 34.755 38.760 34.985 39.065 ;
        RECT 34.235 38.695 34.985 38.760 ;
        RECT 33.205 38.465 34.985 38.695 ;
        RECT 33.205 38.090 33.435 38.465 ;
        RECT 34.235 38.400 34.985 38.465 ;
        RECT 34.755 38.090 34.985 38.400 ;
        RECT 33.205 37.755 34.985 38.090 ;
        RECT 33.205 36.805 33.435 37.755 ;
        RECT 33.655 37.405 33.955 37.470 ;
        RECT 33.595 37.175 34.595 37.405 ;
        RECT 33.655 37.110 33.955 37.175 ;
        RECT 34.755 36.805 34.985 37.755 ;
        RECT 33.205 36.470 34.985 36.805 ;
        RECT 33.205 36.115 33.435 36.470 ;
        RECT 34.755 36.180 34.985 36.470 ;
        RECT 34.235 36.115 34.985 36.180 ;
        RECT 33.205 35.885 34.985 36.115 ;
        RECT 33.205 35.505 33.435 35.885 ;
        RECT 34.235 35.820 34.985 35.885 ;
        RECT 34.755 35.505 34.985 35.820 ;
        RECT 33.205 35.170 34.985 35.505 ;
        RECT 33.205 34.875 33.435 35.170 ;
        RECT 33.655 34.825 33.955 34.890 ;
        RECT 34.755 34.875 34.985 35.170 ;
        RECT 37.095 39.165 37.325 43.575 ;
        RECT 37.590 43.340 38.290 43.435 ;
        RECT 38.735 43.390 38.965 43.575 ;
        RECT 37.530 43.110 38.530 43.340 ;
        RECT 37.590 43.015 38.290 43.110 ;
        RECT 39.225 42.445 39.960 47.495 ;
        RECT 40.290 42.440 41.090 52.455 ;
        RECT 90.140 51.525 91.140 53.535 ;
        RECT 90.140 46.370 90.570 51.525 ;
        RECT 92.025 51.325 108.220 53.535 ;
        RECT 109.135 53.270 109.365 53.330 ;
        RECT 109.065 51.590 109.435 53.270 ;
        RECT 109.135 51.530 109.365 51.590 ;
        RECT 110.335 51.325 126.530 53.535 ;
        RECT 127.355 51.535 128.365 53.335 ;
        RECT 127.425 51.530 127.655 51.535 ;
        RECT 91.125 51.095 109.085 51.325 ;
        RECT 109.415 51.095 127.375 51.325 ;
        RECT 90.710 49.085 91.140 50.890 ;
        RECT 92.025 48.885 108.220 51.095 ;
        RECT 109.135 50.830 109.365 50.890 ;
        RECT 109.065 49.150 109.435 50.830 ;
        RECT 109.135 49.090 109.365 49.150 ;
        RECT 110.335 48.885 126.530 51.095 ;
        RECT 127.365 48.885 127.795 50.890 ;
        RECT 91.125 48.655 127.795 48.885 ;
        RECT 127.935 47.295 128.365 51.535 ;
        RECT 90.710 47.290 129.505 47.295 ;
        RECT 132.440 47.290 133.440 47.295 ;
        RECT 90.710 46.795 133.440 47.290 ;
        RECT 129.430 46.790 133.440 46.795 ;
        RECT 132.440 46.490 133.440 46.790 ;
        RECT 90.140 45.870 127.845 46.370 ;
        RECT 97.175 44.130 109.135 44.360 ;
        RECT 109.465 44.130 121.425 44.360 ;
        RECT 96.895 43.910 97.125 43.970 ;
        RECT 37.855 39.695 38.470 39.760 ;
        RECT 37.530 39.465 38.530 39.695 ;
        RECT 37.855 39.400 38.470 39.465 ;
        RECT 38.735 39.165 38.965 39.415 ;
        RECT 37.095 37.770 38.965 39.165 ;
        RECT 33.595 34.595 34.595 34.825 ;
        RECT 33.205 34.245 33.435 34.545 ;
        RECT 33.655 34.530 33.955 34.595 ;
        RECT 34.755 34.245 34.985 34.545 ;
        RECT 33.205 33.910 34.985 34.245 ;
        RECT 33.205 32.975 33.435 33.910 ;
        RECT 33.655 33.535 33.955 33.600 ;
        RECT 33.595 33.305 34.595 33.535 ;
        RECT 33.655 33.240 33.955 33.305 ;
        RECT 34.755 32.975 34.985 33.910 ;
        RECT 33.205 32.640 34.985 32.975 ;
        RECT 33.205 32.245 33.435 32.640 ;
        RECT 34.755 32.310 34.985 32.640 ;
        RECT 34.235 32.245 34.985 32.310 ;
        RECT 33.205 32.015 34.985 32.245 ;
        RECT 33.205 31.670 33.435 32.015 ;
        RECT 34.235 31.950 34.985 32.015 ;
        RECT 34.755 31.670 34.985 31.950 ;
        RECT 33.205 31.335 34.985 31.670 ;
        RECT 33.205 30.405 33.435 31.335 ;
        RECT 33.655 30.955 33.955 31.020 ;
        RECT 33.595 30.725 34.595 30.955 ;
        RECT 33.655 30.660 33.955 30.725 ;
        RECT 34.755 30.405 34.985 31.335 ;
        RECT 33.205 30.070 34.985 30.405 ;
        RECT 33.205 29.665 33.435 30.070 ;
        RECT 34.755 29.730 34.985 30.070 ;
        RECT 34.235 29.665 34.985 29.730 ;
        RECT 33.205 29.435 34.985 29.665 ;
        RECT 33.205 29.095 33.435 29.435 ;
        RECT 34.235 29.370 34.985 29.435 ;
        RECT 34.755 29.095 34.985 29.370 ;
        RECT 33.205 28.760 34.985 29.095 ;
        RECT 33.205 28.425 33.435 28.760 ;
        RECT 33.655 28.375 33.955 28.440 ;
        RECT 34.755 28.425 34.985 28.760 ;
        RECT 37.095 32.675 37.325 37.770 ;
        RECT 37.590 37.405 38.155 37.470 ;
        RECT 38.735 37.455 38.965 37.770 ;
        RECT 37.530 37.175 38.530 37.405 ;
        RECT 37.590 37.110 38.155 37.175 ;
        RECT 37.855 33.245 38.470 33.310 ;
        RECT 37.530 33.015 38.530 33.245 ;
        RECT 37.855 32.950 38.470 33.015 ;
        RECT 38.735 32.675 38.965 32.965 ;
        RECT 37.095 31.280 38.965 32.675 ;
        RECT 33.595 28.145 34.595 28.375 ;
        RECT 33.205 27.805 33.435 28.095 ;
        RECT 33.655 28.080 33.955 28.145 ;
        RECT 34.755 27.805 34.985 28.095 ;
        RECT 33.205 27.470 34.985 27.805 ;
        RECT 33.205 26.520 33.435 27.470 ;
        RECT 33.655 27.085 33.955 27.150 ;
        RECT 33.595 26.855 34.595 27.085 ;
        RECT 33.655 26.790 33.955 26.855 ;
        RECT 34.755 26.520 34.985 27.470 ;
        RECT 33.205 26.185 34.985 26.520 ;
        RECT 33.205 25.795 33.435 26.185 ;
        RECT 34.755 25.860 34.985 26.185 ;
        RECT 34.235 25.795 34.985 25.860 ;
        RECT 33.205 25.565 34.985 25.795 ;
        RECT 33.205 25.215 33.435 25.565 ;
        RECT 34.235 25.500 34.985 25.565 ;
        RECT 34.755 25.215 34.985 25.500 ;
        RECT 33.205 24.880 34.985 25.215 ;
        RECT 33.205 23.920 33.435 24.880 ;
        RECT 33.655 24.505 33.955 24.570 ;
        RECT 33.595 24.275 34.595 24.505 ;
        RECT 33.655 24.210 33.955 24.275 ;
        RECT 34.755 23.920 34.985 24.880 ;
        RECT 33.205 23.585 34.985 23.920 ;
        RECT 33.205 23.215 33.435 23.585 ;
        RECT 34.755 23.280 34.985 23.585 ;
        RECT 34.235 23.215 34.985 23.280 ;
        RECT 33.205 22.985 34.985 23.215 ;
        RECT 33.205 22.670 33.435 22.985 ;
        RECT 34.235 22.920 34.985 22.985 ;
        RECT 34.755 22.670 34.985 22.920 ;
        RECT 33.205 22.335 34.985 22.670 ;
        RECT 33.205 21.975 33.435 22.335 ;
        RECT 33.655 21.925 33.955 21.990 ;
        RECT 34.755 21.975 34.985 22.335 ;
        RECT 37.095 26.270 37.325 31.280 ;
        RECT 37.590 30.955 38.155 31.020 ;
        RECT 38.735 31.005 38.965 31.280 ;
        RECT 37.530 30.725 38.530 30.955 ;
        RECT 37.590 30.660 38.155 30.725 ;
        RECT 37.855 26.795 38.470 26.860 ;
        RECT 37.530 26.565 38.530 26.795 ;
        RECT 37.855 26.500 38.470 26.565 ;
        RECT 38.735 26.270 38.965 26.515 ;
        RECT 37.095 24.875 38.965 26.270 ;
        RECT 33.595 21.695 34.595 21.925 ;
        RECT 33.205 21.370 33.435 21.645 ;
        RECT 33.655 21.630 33.955 21.695 ;
        RECT 34.755 21.370 34.985 21.645 ;
        RECT 33.205 21.035 34.985 21.370 ;
        RECT 33.205 20.060 33.435 21.035 ;
        RECT 33.655 20.635 33.955 20.700 ;
        RECT 33.595 20.405 34.595 20.635 ;
        RECT 33.655 20.340 33.955 20.405 ;
        RECT 34.755 20.060 34.985 21.035 ;
        RECT 33.205 19.725 34.985 20.060 ;
        RECT 33.205 19.345 33.435 19.725 ;
        RECT 34.755 19.410 34.985 19.725 ;
        RECT 34.235 19.345 34.985 19.410 ;
        RECT 33.205 19.115 34.985 19.345 ;
        RECT 33.205 18.760 33.435 19.115 ;
        RECT 34.235 19.050 34.985 19.115 ;
        RECT 34.755 18.760 34.985 19.050 ;
        RECT 33.205 18.425 34.985 18.760 ;
        RECT 33.205 17.465 33.435 18.425 ;
        RECT 33.655 18.055 33.955 18.120 ;
        RECT 33.595 17.825 34.595 18.055 ;
        RECT 33.655 17.760 33.955 17.825 ;
        RECT 34.755 17.465 34.985 18.425 ;
        RECT 33.205 17.130 34.985 17.465 ;
        RECT 33.205 16.765 33.435 17.130 ;
        RECT 34.755 16.830 34.985 17.130 ;
        RECT 34.235 16.765 34.985 16.830 ;
        RECT 33.205 16.535 34.985 16.765 ;
        RECT 33.205 16.130 33.435 16.535 ;
        RECT 34.235 16.470 34.985 16.535 ;
        RECT 34.755 16.130 34.985 16.470 ;
        RECT 33.205 15.795 34.985 16.130 ;
        RECT 33.205 15.525 33.435 15.795 ;
        RECT 33.655 15.475 33.955 15.540 ;
        RECT 34.235 15.475 34.535 15.540 ;
        RECT 34.755 15.525 34.985 15.795 ;
        RECT 37.095 19.720 37.325 24.875 ;
        RECT 37.590 24.505 38.155 24.570 ;
        RECT 38.735 24.555 38.965 24.875 ;
        RECT 37.530 24.275 38.530 24.505 ;
        RECT 37.590 24.210 38.155 24.275 ;
        RECT 39.795 21.300 40.550 39.760 ;
        RECT 96.655 38.240 97.185 43.910 ;
        RECT 96.895 37.970 97.125 38.240 ;
        RECT 100.415 37.840 105.840 44.130 ;
        RECT 109.185 39.785 109.415 43.970 ;
        RECT 109.125 38.190 109.485 39.785 ;
        RECT 109.185 37.970 109.415 38.190 ;
        RECT 112.935 37.840 118.370 44.130 ;
        RECT 121.475 43.910 121.705 43.970 ;
        RECT 121.415 38.305 121.945 43.910 ;
        RECT 121.475 37.970 121.705 38.305 ;
        RECT 97.205 37.810 109.125 37.840 ;
        RECT 109.475 37.810 121.415 37.840 ;
        RECT 97.175 37.580 109.135 37.810 ;
        RECT 109.465 37.580 121.425 37.810 ;
        RECT 97.205 37.555 109.125 37.580 ;
        RECT 109.475 37.555 121.415 37.580 ;
        RECT 97.255 36.875 110.570 37.270 ;
        RECT 90.240 36.375 93.220 36.430 ;
        RECT 90.230 36.145 93.230 36.375 ;
        RECT 89.840 35.100 90.070 36.095 ;
        RECT 93.390 35.190 93.685 36.095 ;
        RECT 108.020 35.340 121.365 35.785 ;
        RECT 93.330 35.100 93.690 35.190 ;
        RECT 89.840 32.115 93.690 35.100 ;
        RECT 97.180 34.985 109.120 35.015 ;
        RECT 109.470 34.985 121.410 35.010 ;
        RECT 97.170 34.755 109.130 34.985 ;
        RECT 109.460 34.755 121.420 34.985 ;
        RECT 97.180 34.730 109.120 34.755 ;
        RECT 96.890 34.535 97.120 34.595 ;
        RECT 89.840 31.135 90.070 32.115 ;
        RECT 93.330 31.195 93.690 32.115 ;
        RECT 93.390 31.135 93.685 31.195 ;
        RECT 90.230 30.855 93.230 31.085 ;
        RECT 96.125 28.830 97.180 34.535 ;
        RECT 96.890 28.595 97.120 28.830 ;
        RECT 100.390 28.440 105.825 34.730 ;
        RECT 109.470 34.725 121.410 34.755 ;
        RECT 109.180 34.380 109.410 34.595 ;
        RECT 109.120 32.785 109.480 34.380 ;
        RECT 109.180 28.595 109.410 32.785 ;
        RECT 89.100 27.835 91.985 28.365 ;
        RECT 97.170 28.180 109.130 28.440 ;
        RECT 109.470 28.435 111.970 28.445 ;
        RECT 112.890 28.435 118.325 34.725 ;
        RECT 121.470 34.535 121.700 34.595 ;
        RECT 121.405 29.175 122.265 34.535 ;
        RECT 121.470 28.595 121.700 29.175 ;
        RECT 109.460 28.205 121.420 28.435 ;
        RECT 109.470 28.185 111.970 28.205 ;
        RECT 89.110 26.685 123.900 27.190 ;
        RECT 39.775 21.010 40.570 21.300 ;
        RECT 37.850 20.345 38.470 20.410 ;
        RECT 37.530 20.115 38.530 20.345 ;
        RECT 37.850 20.050 38.470 20.115 ;
        RECT 38.735 19.720 38.965 20.065 ;
        RECT 37.095 18.325 38.965 19.720 ;
        RECT 37.095 16.840 37.325 18.325 ;
        RECT 37.590 18.055 38.205 18.120 ;
        RECT 38.735 18.105 38.965 18.325 ;
        RECT 37.530 17.825 38.530 18.055 ;
        RECT 37.590 17.760 38.205 17.825 ;
        RECT 37.855 17.440 38.470 17.505 ;
        RECT 37.530 17.210 38.530 17.440 ;
        RECT 37.855 17.145 38.470 17.210 ;
        RECT 38.735 16.840 38.965 17.160 ;
        RECT 33.595 15.245 34.595 15.475 ;
        RECT 37.095 15.445 38.965 16.840 ;
        RECT 33.655 15.180 33.955 15.245 ;
        RECT 34.235 15.180 34.535 15.245 ;
        RECT 37.095 15.175 37.325 15.445 ;
        RECT 37.590 15.150 38.205 15.215 ;
        RECT 38.735 15.200 38.965 15.445 ;
        RECT 37.530 14.920 38.530 15.150 ;
        RECT 37.590 14.855 38.205 14.920 ;
        RECT 39.795 14.615 40.550 21.010 ;
      LAYER met2 ;
        RECT 85.860 148.285 99.265 149.400 ;
        RECT 85.860 148.280 87.130 148.285 ;
        RECT 80.160 140.250 83.635 142.365 ;
        RECT 86.305 140.250 87.130 148.280 ;
        RECT 90.090 146.420 103.495 146.920 ;
        RECT 90.090 143.820 90.450 146.420 ;
        RECT 94.470 143.820 94.830 146.420 ;
        RECT 80.160 140.245 87.130 140.250 ;
        RECT 43.285 138.245 87.130 140.245 ;
        RECT 45.315 130.530 45.745 134.110 ;
        RECT 63.770 132.320 64.040 138.245 ;
        RECT 45.315 130.010 46.910 130.530 ;
        RECT 49.405 130.015 51.210 130.515 ;
        RECT 74.725 130.015 76.550 130.515 ;
        RECT 44.945 119.325 47.825 119.750 ;
        RECT 48.035 118.455 48.295 118.460 ;
        RECT 48.020 114.365 48.310 118.455 ;
        RECT 50.780 117.805 51.210 130.015 ;
        RECT 51.360 129.090 53.290 129.590 ;
        RECT 51.360 124.240 51.790 129.090 ;
        RECT 76.120 124.240 76.550 130.015 ;
        RECT 82.070 129.590 82.500 134.110 ;
        RECT 86.305 131.245 87.130 138.245 ;
        RECT 92.300 138.125 92.620 143.225 ;
        RECT 87.915 131.940 88.235 137.040 ;
        RECT 96.680 131.940 97.000 137.040 ;
        RECT 88.305 131.430 89.705 131.790 ;
        RECT 90.495 131.430 91.895 131.790 ;
        RECT 92.685 131.430 94.085 131.790 ;
        RECT 94.875 131.430 96.275 131.790 ;
        RECT 88.305 129.965 88.805 131.430 ;
        RECT 76.700 129.090 78.570 129.590 ;
        RECT 80.395 129.090 82.500 129.590 ;
        RECT 63.810 121.310 64.090 123.120 ;
        RECT 51.910 120.135 52.960 121.110 ;
        RECT 62.675 117.900 63.725 118.945 ;
        RECT 64.175 117.895 65.225 120.550 ;
        RECT 74.970 118.570 76.020 121.110 ;
        RECT 76.700 117.805 77.130 129.090 ;
        RECT 89.545 127.545 90.045 129.020 ;
        RECT 90.495 128.420 90.995 131.430 ;
        RECT 91.735 127.545 92.235 130.565 ;
        RECT 92.685 128.420 93.185 131.430 ;
        RECT 93.925 127.545 94.425 130.565 ;
        RECT 94.875 129.965 95.375 131.430 ;
        RECT 96.115 127.545 96.615 129.020 ;
        RECT 50.780 114.935 51.785 117.805 ;
        RECT 63.805 115.905 64.095 117.700 ;
        RECT 50.780 112.050 51.795 114.935 ;
        RECT 76.110 112.345 77.130 117.805 ;
        RECT 86.390 114.295 87.130 127.255 ;
        RECT 88.645 127.185 90.045 127.545 ;
        RECT 90.835 127.185 92.235 127.545 ;
        RECT 93.025 127.185 94.425 127.545 ;
        RECT 95.215 127.185 96.615 127.545 ;
        RECT 87.920 121.935 88.240 127.035 ;
        RECT 96.680 121.935 97.000 127.035 ;
        RECT 92.300 116.135 92.620 121.235 ;
        RECT 102.995 119.265 103.495 146.420 ;
        RECT 103.950 129.965 105.410 130.565 ;
        RECT 121.325 121.830 130.975 121.845 ;
        RECT 104.680 120.285 130.975 121.830 ;
        RECT 104.680 120.275 122.995 120.285 ;
        RECT 102.995 118.765 120.715 119.265 ;
        RECT 90.090 115.155 97.090 115.160 ;
        RECT 102.995 115.155 103.495 118.765 ;
        RECT 90.090 114.660 103.495 115.155 ;
        RECT 38.295 111.885 39.480 111.935 ;
        RECT 38.295 110.430 47.185 111.885 ;
        RECT 51.885 111.335 54.285 111.725 ;
        RECT 64.175 111.345 66.575 111.735 ;
        RECT 85.675 111.210 87.160 114.295 ;
        RECT 90.090 112.055 90.450 114.660 ;
        RECT 94.465 112.055 94.825 114.660 ;
        RECT 96.450 114.655 103.495 114.660 ;
        RECT 112.095 114.165 112.355 118.765 ;
        RECT 114.185 111.595 114.445 117.385 ;
        RECT 116.275 114.165 116.535 118.765 ;
        RECT 118.365 111.595 118.625 117.385 ;
        RECT 120.455 114.165 120.715 118.765 ;
        RECT 121.560 112.695 122.995 120.275 ;
        RECT 125.880 114.165 126.310 120.010 ;
        RECT 126.815 118.470 127.135 119.170 ;
        RECT 126.810 114.090 127.130 114.790 ;
        RECT 127.695 113.345 128.090 119.990 ;
        RECT 121.495 111.770 129.555 112.165 ;
        RECT 38.295 109.885 78.495 110.430 ;
        RECT 85.675 110.390 99.210 111.210 ;
        RECT 85.675 110.360 87.160 110.390 ;
        RECT 110.730 110.315 121.045 111.595 ;
        RECT 38.295 109.880 44.065 109.885 ;
        RECT 38.295 109.830 39.480 109.880 ;
        RECT 74.665 108.790 78.495 109.885 ;
        RECT 86.665 108.790 87.400 108.800 ;
        RECT 74.665 108.760 87.400 108.790 ;
        RECT 74.665 108.755 88.045 108.760 ;
        RECT 47.970 108.630 48.870 108.685 ;
        RECT 47.970 108.130 70.335 108.630 ;
        RECT 47.970 108.080 48.870 108.130 ;
        RECT 69.835 94.185 70.335 108.130 ;
        RECT 74.665 108.140 126.120 108.755 ;
        RECT 74.665 106.045 87.400 108.140 ;
        RECT 87.970 106.305 88.290 106.905 ;
        RECT 97.690 106.305 97.950 108.140 ;
        RECT 117.070 106.305 117.330 108.140 ;
        RECT 126.730 106.305 127.050 106.905 ;
        RECT 74.665 105.995 77.985 106.045 ;
        RECT 86.665 102.290 87.400 106.045 ;
        RECT 107.350 105.425 107.670 106.025 ;
        RECT 107.350 104.255 107.670 104.855 ;
        RECT 87.970 103.375 88.290 103.975 ;
        RECT 86.335 102.285 87.870 102.290 ;
        RECT 97.690 102.285 97.950 103.975 ;
        RECT 117.070 102.285 117.330 103.975 ;
        RECT 126.730 103.375 127.050 103.975 ;
        RECT 86.335 101.200 126.260 102.285 ;
        RECT 129.160 100.165 129.555 111.770 ;
        RECT 80.635 99.130 83.475 99.830 ;
        RECT 128.725 99.565 129.555 100.165 ;
        RECT 80.635 98.290 83.505 99.130 ;
        RECT 118.410 98.800 119.520 98.850 ;
        RECT 80.330 98.260 87.100 98.290 ;
        RECT 107.670 98.260 119.520 98.800 ;
        RECT 80.330 97.465 119.520 98.260 ;
        RECT 80.330 97.435 87.100 97.465 ;
        RECT 69.835 94.085 79.845 94.185 ;
        RECT 80.570 94.085 80.830 95.945 ;
        RECT 82.860 95.495 83.120 97.435 ;
        RECT 69.835 93.840 81.155 94.085 ;
        RECT 69.835 93.685 79.845 93.840 ;
        RECT 80.895 91.695 81.155 93.840 ;
        RECT 83.475 92.275 83.735 95.940 ;
        RECT 85.765 95.490 86.025 97.435 ;
        RECT 89.925 92.275 90.185 95.895 ;
        RECT 92.215 95.495 92.475 97.465 ;
        RECT 96.375 92.275 96.635 95.895 ;
        RECT 98.665 95.495 98.925 97.465 ;
        RECT 102.825 92.275 103.085 95.895 ;
        RECT 105.115 95.495 105.375 97.465 ;
        RECT 107.675 96.905 119.520 97.465 ;
        RECT 107.675 96.895 112.605 96.905 ;
        RECT 108.235 95.230 108.555 96.030 ;
        RECT 109.555 95.410 109.815 96.895 ;
        RECT 110.815 95.230 111.135 96.030 ;
        RECT 114.180 95.230 114.440 96.905 ;
        RECT 115.480 96.810 115.740 96.905 ;
        RECT 118.410 96.855 119.520 96.905 ;
        RECT 112.275 94.630 114.070 95.055 ;
        RECT 114.545 94.630 116.340 95.055 ;
        RECT 111.115 92.450 117.085 93.400 ;
        RECT 82.185 91.875 85.025 92.275 ;
        RECT 88.635 91.875 91.475 92.275 ;
        RECT 95.085 91.875 97.925 92.275 ;
        RECT 101.535 91.875 104.375 92.275 ;
        RECT 98.925 91.695 99.245 91.715 ;
        RECT 80.895 91.295 86.315 91.695 ;
        RECT 87.345 91.295 92.765 91.695 ;
        RECT 93.795 91.295 99.245 91.695 ;
        RECT 100.245 91.295 105.665 91.695 ;
        RECT 106.695 91.295 109.185 91.695 ;
        RECT 74.665 90.550 77.980 90.600 ;
        RECT 74.665 89.495 107.980 90.550 ;
        RECT 74.665 89.485 81.165 89.495 ;
        RECT 74.665 89.435 77.980 89.485 ;
        RECT 108.785 87.685 109.185 91.295 ;
        RECT 111.115 86.445 111.885 92.450 ;
        RECT 112.740 88.715 113.110 91.815 ;
        RECT 116.280 89.640 117.085 92.450 ;
        RECT 151.810 88.235 152.710 103.925 ;
        RECT 151.790 87.385 152.730 88.235 ;
        RECT 151.810 87.360 152.710 87.385 ;
        RECT 113.645 86.445 116.305 87.170 ;
        RECT 84.535 86.055 116.305 86.445 ;
        RECT 84.535 85.785 117.190 86.055 ;
        RECT 84.920 83.490 85.180 85.785 ;
        RECT 87.490 83.490 87.770 84.590 ;
        RECT 90.070 83.490 90.350 84.590 ;
        RECT 92.660 83.490 92.920 85.785 ;
        RECT 95.230 83.490 95.510 84.590 ;
        RECT 97.810 83.490 98.090 84.590 ;
        RECT 100.400 83.490 100.660 85.785 ;
        RECT 102.970 83.490 103.250 84.590 ;
        RECT 105.550 83.490 105.830 84.590 ;
        RECT 108.140 83.490 108.400 85.785 ;
        RECT 110.710 83.490 110.990 84.590 ;
        RECT 113.290 83.485 113.570 84.585 ;
        RECT 115.880 83.490 116.140 85.785 ;
        RECT 93.315 82.715 93.575 82.725 ;
        RECT 99.795 82.715 100.055 82.725 ;
        RECT 115.205 82.715 115.465 82.725 ;
        RECT 83.520 82.115 115.585 82.715 ;
        RECT 83.520 75.565 84.120 82.115 ;
        RECT 85.580 82.105 85.840 82.115 ;
        RECT 99.110 82.110 99.370 82.115 ;
        RECT 107.535 82.105 107.795 82.115 ;
        RECT 108.815 82.110 109.075 82.115 ;
        RECT 88.760 80.610 89.080 81.710 ;
        RECT 96.500 80.610 96.820 81.710 ;
        RECT 104.240 80.610 104.560 81.710 ;
        RECT 111.980 80.610 112.300 81.710 ;
        RECT 85.275 80.145 85.775 80.505 ;
        RECT 86.565 80.145 87.485 80.505 ;
        RECT 91.725 80.145 92.225 80.505 ;
        RECT 94.305 80.145 95.225 80.505 ;
        RECT 99.465 80.145 99.965 80.505 ;
        RECT 102.045 80.145 102.965 80.505 ;
        RECT 107.205 80.145 107.705 80.505 ;
        RECT 109.785 80.145 110.785 80.505 ;
        RECT 114.945 80.145 115.445 80.505 ;
        RECT 85.275 79.505 85.535 80.145 ;
        RECT 85.035 79.145 85.535 79.505 ;
        RECT 86.565 78.780 86.825 80.145 ;
        RECT 91.725 79.505 91.985 80.145 ;
        RECT 87.615 79.145 88.115 79.505 ;
        RECT 91.485 79.145 91.985 79.505 ;
        RECT 85.035 78.420 85.535 78.780 ;
        RECT 86.325 78.420 86.825 78.780 ;
        RECT 85.275 77.650 85.535 78.420 ;
        RECT 87.855 77.650 88.115 79.145 ;
        RECT 94.305 78.780 94.565 80.145 ;
        RECT 99.465 79.505 99.725 80.145 ;
        RECT 95.355 79.145 95.855 79.505 ;
        RECT 99.225 79.145 99.725 79.505 ;
        RECT 90.195 78.420 90.695 78.780 ;
        RECT 94.065 78.420 94.565 78.780 ;
        RECT 90.435 77.650 90.695 78.420 ;
        RECT 95.595 77.650 95.855 79.145 ;
        RECT 102.045 78.780 102.305 80.145 ;
        RECT 107.205 79.505 107.465 80.145 ;
        RECT 103.095 79.145 103.595 79.505 ;
        RECT 106.965 79.145 107.465 79.505 ;
        RECT 97.935 78.420 98.435 78.780 ;
        RECT 101.805 78.420 102.305 78.780 ;
        RECT 98.175 77.650 98.435 78.420 ;
        RECT 103.335 77.650 103.595 79.145 ;
        RECT 109.785 78.780 110.045 80.145 ;
        RECT 114.945 79.505 115.205 80.145 ;
        RECT 110.835 79.145 111.335 79.505 ;
        RECT 114.705 79.145 115.205 79.505 ;
        RECT 105.675 78.420 106.175 78.780 ;
        RECT 109.545 78.420 110.045 78.780 ;
        RECT 105.915 77.650 106.175 78.420 ;
        RECT 111.075 77.650 111.335 79.145 ;
        RECT 113.415 78.420 113.915 78.780 ;
        RECT 113.655 77.650 113.915 78.420 ;
        RECT 85.275 77.290 85.775 77.650 ;
        RECT 87.855 77.290 88.355 77.650 ;
        RECT 90.435 77.290 91.060 77.650 ;
        RECT 95.595 77.290 96.095 77.650 ;
        RECT 98.175 77.290 98.805 77.650 ;
        RECT 103.335 77.290 103.835 77.650 ;
        RECT 105.915 77.290 106.575 77.650 ;
        RECT 111.075 77.290 111.575 77.650 ;
        RECT 113.655 77.290 114.155 77.650 ;
        RECT 86.200 76.085 86.480 77.185 ;
        RECT 91.360 76.085 91.640 77.185 ;
        RECT 93.940 76.085 94.220 77.185 ;
        RECT 99.100 76.085 99.380 77.185 ;
        RECT 101.680 76.085 101.960 77.185 ;
        RECT 106.840 76.085 107.120 77.185 ;
        RECT 109.420 76.085 109.700 77.185 ;
        RECT 114.580 76.085 114.860 77.185 ;
        RECT 97.170 75.565 97.430 75.575 ;
        RECT 103.635 75.565 103.895 75.570 ;
        RECT 83.520 74.965 113.560 75.565 ;
        RECT 88.145 74.960 88.405 74.965 ;
        RECT 89.455 74.950 89.715 74.965 ;
        RECT 95.910 74.960 96.170 74.965 ;
        RECT 104.945 74.960 105.205 74.965 ;
        RECT 84.890 73.205 85.210 74.305 ;
        RECT 74.665 72.060 77.985 72.115 ;
        RECT 74.665 72.050 84.930 72.060 ;
        RECT 88.790 72.050 89.050 74.305 ;
        RECT 92.630 73.205 92.950 74.305 ;
        RECT 96.535 72.050 96.795 74.305 ;
        RECT 100.370 73.205 100.690 74.305 ;
        RECT 104.270 72.050 104.530 74.305 ;
        RECT 108.110 73.205 108.430 74.305 ;
        RECT 112.010 72.050 112.270 74.305 ;
        RECT 115.850 73.205 116.170 74.305 ;
        RECT 116.920 72.050 117.190 85.785 ;
        RECT 74.665 71.080 117.765 72.050 ;
        RECT 74.665 71.030 77.985 71.080 ;
        RECT 69.815 61.365 70.840 61.415 ;
        RECT 39.225 59.460 70.840 61.365 ;
        RECT 9.515 52.100 11.515 52.150 ;
        RECT 13.390 52.100 14.360 52.795 ;
        RECT 39.225 52.400 41.130 59.460 ;
        RECT 69.815 59.410 70.840 59.460 ;
        RECT 129.510 57.025 130.680 57.070 ;
        RECT 88.630 55.025 130.680 57.025 ;
        RECT 9.515 52.020 14.360 52.100 ;
        RECT 9.515 51.750 28.365 52.020 ;
        RECT 9.515 50.100 14.360 51.750 ;
        RECT 28.095 51.135 28.365 51.750 ;
        RECT 15.515 50.680 16.615 51.000 ;
        RECT 28.095 50.970 29.480 51.135 ;
        RECT 31.950 51.110 35.710 51.915 ;
        RECT 39.215 51.900 41.130 52.400 ;
        RECT 25.800 50.710 29.480 50.970 ;
        RECT 24.425 50.295 25.025 50.415 ;
        RECT 9.515 50.050 11.515 50.100 ;
        RECT 13.390 47.100 14.360 50.100 ;
        RECT 22.455 50.035 22.815 50.275 ;
        RECT 21.455 49.775 22.815 50.035 ;
        RECT 24.425 50.035 25.035 50.295 ;
        RECT 18.395 49.410 19.495 49.690 ;
        RECT 21.455 49.535 21.815 49.775 ;
        RECT 19.600 48.745 19.960 48.985 ;
        RECT 19.600 48.485 21.090 48.745 ;
        RECT 13.390 46.840 16.615 47.100 ;
        RECT 13.390 39.360 14.360 46.840 ;
        RECT 15.515 42.940 16.615 43.260 ;
        RECT 17.275 40.035 17.875 48.390 ;
        RECT 20.730 48.245 21.090 48.485 ;
        RECT 22.920 46.810 24.020 47.130 ;
        RECT 19.600 46.165 19.960 46.405 ;
        RECT 19.600 45.905 21.815 46.165 ;
        RECT 21.455 45.665 21.815 45.905 ;
        RECT 22.455 44.875 22.815 45.615 ;
        RECT 20.730 44.615 22.815 44.875 ;
        RECT 18.395 44.250 19.495 44.530 ;
        RECT 20.730 44.375 21.090 44.615 ;
        RECT 24.425 43.905 25.025 50.035 ;
        RECT 28.095 48.475 29.480 50.710 ;
        RECT 25.795 48.120 26.895 48.400 ;
        RECT 28.095 46.715 28.755 48.475 ;
        RECT 31.025 47.570 34.125 47.940 ;
        RECT 34.760 46.715 35.710 51.110 ;
        RECT 36.940 49.375 37.365 51.170 ;
        RECT 39.215 50.570 41.110 51.900 ;
        RECT 39.120 50.310 41.110 50.570 ;
        RECT 39.215 49.270 41.110 50.310 ;
        RECT 37.540 49.010 41.110 49.270 ;
        RECT 36.940 47.105 37.365 48.900 ;
        RECT 39.215 47.435 41.110 49.010 ;
        RECT 28.095 45.945 35.710 46.715 ;
        RECT 25.800 45.540 26.900 45.820 ;
        RECT 24.420 43.645 25.025 43.905 ;
        RECT 24.425 42.625 25.025 43.645 ;
        RECT 28.095 43.230 28.755 45.945 ;
        RECT 37.540 45.645 38.340 45.965 ;
        RECT 39.205 44.645 41.110 47.435 ;
        RECT 90.660 47.310 91.090 50.890 ;
        RECT 109.115 49.100 109.385 55.025 ;
        RECT 129.510 54.970 130.680 55.025 ;
        RECT 90.660 46.790 92.255 47.310 ;
        RECT 94.750 46.795 96.555 47.295 ;
        RECT 120.070 46.795 121.895 47.295 ;
        RECT 37.720 44.385 41.110 44.645 ;
        RECT 29.935 43.330 34.005 43.730 ;
        RECT 25.800 42.970 28.755 43.230 ;
        RECT 22.455 42.295 22.815 42.535 ;
        RECT 24.415 42.365 25.025 42.625 ;
        RECT 21.455 42.035 22.815 42.295 ;
        RECT 18.395 41.670 19.495 41.950 ;
        RECT 21.455 41.795 21.815 42.035 ;
        RECT 19.600 41.005 19.960 41.405 ;
        RECT 19.600 40.745 21.090 41.005 ;
        RECT 20.730 40.505 21.090 40.745 ;
        RECT 17.270 39.775 17.875 40.035 ;
        RECT 13.390 39.100 16.615 39.360 ;
        RECT 13.390 31.625 14.360 39.100 ;
        RECT 17.275 38.725 17.875 39.775 ;
        RECT 22.920 39.070 24.020 39.390 ;
        RECT 17.275 38.465 17.880 38.725 ;
        RECT 15.515 35.200 16.615 35.520 ;
        RECT 17.275 32.260 17.875 38.465 ;
        RECT 19.600 38.425 19.960 38.665 ;
        RECT 19.600 38.165 21.815 38.425 ;
        RECT 21.455 37.925 21.815 38.165 ;
        RECT 22.455 37.135 22.815 37.795 ;
        RECT 20.730 36.875 22.815 37.135 ;
        RECT 18.395 36.510 19.495 36.790 ;
        RECT 20.730 36.635 21.090 36.875 ;
        RECT 24.425 34.885 25.025 42.365 ;
        RECT 25.800 40.380 26.900 40.660 ;
        RECT 25.800 37.800 26.900 38.080 ;
        RECT 28.095 35.490 28.755 42.970 ;
        RECT 25.800 35.230 28.755 35.490 ;
        RECT 22.455 34.555 22.815 34.795 ;
        RECT 21.455 34.295 22.815 34.555 ;
        RECT 24.425 34.625 25.035 34.885 ;
        RECT 18.395 33.930 19.495 34.210 ;
        RECT 21.455 34.055 21.815 34.295 ;
        RECT 24.425 34.200 25.025 34.625 ;
        RECT 24.420 33.940 25.025 34.200 ;
        RECT 19.600 33.265 19.960 33.635 ;
        RECT 19.600 33.005 21.090 33.265 ;
        RECT 20.730 32.765 21.090 33.005 ;
        RECT 17.275 32.000 17.885 32.260 ;
        RECT 13.390 31.365 16.615 31.625 ;
        RECT 13.390 23.880 14.360 31.365 ;
        RECT 17.275 31.000 17.875 32.000 ;
        RECT 22.920 31.330 24.020 31.650 ;
        RECT 17.270 30.740 17.875 31.000 ;
        RECT 15.515 27.460 16.615 27.780 ;
        RECT 17.275 24.545 17.875 30.740 ;
        RECT 19.600 30.685 19.960 30.925 ;
        RECT 19.600 30.425 21.815 30.685 ;
        RECT 21.455 30.185 21.815 30.425 ;
        RECT 22.455 29.395 22.815 30.055 ;
        RECT 20.730 29.135 22.815 29.395 ;
        RECT 18.395 28.770 19.495 29.050 ;
        RECT 20.730 28.895 21.090 29.135 ;
        RECT 24.425 28.405 25.025 33.940 ;
        RECT 25.800 32.640 26.900 32.920 ;
        RECT 25.800 30.060 26.900 30.340 ;
        RECT 24.425 28.145 25.035 28.405 ;
        RECT 22.455 26.815 22.815 27.055 ;
        RECT 21.455 26.555 22.815 26.815 ;
        RECT 18.395 26.190 19.495 26.470 ;
        RECT 21.455 26.315 21.815 26.555 ;
        RECT 19.600 25.525 19.960 25.890 ;
        RECT 19.600 25.265 21.090 25.525 ;
        RECT 20.730 25.025 21.090 25.265 ;
        RECT 17.260 24.285 17.875 24.545 ;
        RECT 13.390 23.620 16.615 23.880 ;
        RECT 13.390 19.145 14.360 23.620 ;
        RECT 17.275 23.235 17.875 24.285 ;
        RECT 22.920 23.590 24.020 23.910 ;
        RECT 17.270 22.975 17.875 23.235 ;
        RECT 15.515 19.720 16.615 20.040 ;
        RECT 17.275 18.950 17.875 22.975 ;
        RECT 19.600 22.945 19.960 23.185 ;
        RECT 19.600 22.685 21.815 22.945 ;
        RECT 21.455 22.445 21.815 22.685 ;
        RECT 22.455 21.655 22.815 22.315 ;
        RECT 20.730 21.395 22.815 21.655 ;
        RECT 18.395 21.030 19.495 21.310 ;
        RECT 20.730 21.155 21.090 21.395 ;
        RECT 24.425 20.670 25.025 28.145 ;
        RECT 28.095 27.750 28.755 35.230 ;
        RECT 25.800 27.490 28.755 27.750 ;
        RECT 25.800 24.900 26.900 25.180 ;
        RECT 25.800 22.320 26.900 22.600 ;
        RECT 19.600 20.365 19.960 20.605 ;
        RECT 22.455 20.365 22.815 20.605 ;
        RECT 24.415 20.410 25.025 20.670 ;
        RECT 19.600 20.105 21.090 20.365 ;
        RECT 20.730 19.865 21.090 20.105 ;
        RECT 21.455 20.105 22.815 20.365 ;
        RECT 21.455 19.865 21.815 20.105 ;
        RECT 24.425 18.950 25.025 20.410 ;
        RECT 28.095 20.010 28.755 27.490 ;
        RECT 25.800 19.750 28.755 20.010 ;
        RECT 28.095 19.365 28.755 19.750 ;
        RECT 17.275 18.350 25.025 18.950 ;
        RECT 31.805 14.815 32.860 42.315 ;
        RECT 33.605 41.030 34.005 43.330 ;
        RECT 37.540 43.065 38.340 43.385 ;
        RECT 39.205 42.505 41.110 44.385 ;
        RECT 39.770 42.500 41.110 42.505 ;
        RECT 39.770 40.210 40.575 42.500 ;
        RECT 33.605 34.580 34.005 40.000 ;
        RECT 39.775 39.710 40.570 40.210 ;
        RECT 37.805 39.450 40.570 39.710 ;
        RECT 34.185 37.420 34.585 38.710 ;
        RECT 34.185 37.160 38.205 37.420 ;
        RECT 34.185 35.870 34.585 37.160 ;
        RECT 33.605 28.130 34.005 33.550 ;
        RECT 39.775 33.260 40.570 39.450 ;
        RECT 90.290 36.105 93.170 36.530 ;
        RECT 93.380 35.235 93.640 35.240 ;
        RECT 37.805 33.000 40.570 33.260 ;
        RECT 34.185 30.970 34.585 32.260 ;
        RECT 34.185 30.710 38.205 30.970 ;
        RECT 34.185 29.420 34.585 30.710 ;
        RECT 33.605 21.680 34.005 27.100 ;
        RECT 39.775 26.810 40.570 33.000 ;
        RECT 37.805 26.550 40.570 26.810 ;
        RECT 57.505 28.660 59.430 32.815 ;
        RECT 93.365 31.145 93.655 35.235 ;
        RECT 96.125 34.585 96.555 46.795 ;
        RECT 96.705 45.870 98.635 46.370 ;
        RECT 96.705 41.020 97.135 45.870 ;
        RECT 121.465 41.020 121.895 46.795 ;
        RECT 127.415 46.370 127.845 50.890 ;
        RECT 132.490 46.440 133.390 47.345 ;
        RECT 122.045 45.870 123.915 46.370 ;
        RECT 125.740 45.870 127.845 46.370 ;
        RECT 109.155 38.090 109.435 39.900 ;
        RECT 97.255 36.915 98.305 37.890 ;
        RECT 108.020 34.680 109.070 35.725 ;
        RECT 109.520 34.675 110.570 37.330 ;
        RECT 120.315 35.350 121.365 37.890 ;
        RECT 122.045 34.585 122.475 45.870 ;
        RECT 151.810 40.385 152.710 65.190 ;
        RECT 96.125 31.715 97.130 34.585 ;
        RECT 109.150 32.685 109.440 34.480 ;
        RECT 96.125 28.830 97.140 31.715 ;
        RECT 121.455 29.125 122.475 34.585 ;
        RECT 88.620 28.660 92.530 28.665 ;
        RECT 57.505 27.210 92.530 28.660 ;
        RECT 97.230 28.115 99.630 28.505 ;
        RECT 109.520 28.125 111.920 28.515 ;
        RECT 57.505 26.735 123.840 27.210 ;
        RECT 87.235 26.665 123.840 26.735 ;
        RECT 87.235 26.660 88.635 26.665 ;
        RECT 34.185 24.520 34.585 25.810 ;
        RECT 34.185 24.260 38.205 24.520 ;
        RECT 34.185 22.970 34.585 24.260 ;
        RECT 39.775 21.435 40.570 26.550 ;
        RECT 33.605 15.490 34.005 20.650 ;
        RECT 39.745 20.360 40.600 21.435 ;
        RECT 37.800 20.100 40.600 20.360 ;
        RECT 34.185 18.070 34.585 19.360 ;
        RECT 34.185 17.810 38.250 18.070 ;
        RECT 34.185 16.520 34.585 17.810 ;
        RECT 39.745 17.455 40.600 20.100 ;
        RECT 37.805 17.195 40.600 17.455 ;
        RECT 33.605 15.230 36.790 15.490 ;
        RECT 35.890 15.165 36.790 15.230 ;
        RECT 35.890 14.905 38.255 15.165 ;
        RECT 35.890 13.240 36.790 14.905 ;
        RECT 39.745 14.665 40.600 17.195 ;
      LAYER met3 ;
        RECT 87.390 148.440 98.350 149.340 ;
        RECT 80.545 139.270 83.030 141.865 ;
        RECT 92.250 138.605 92.670 143.200 ;
        RECT 92.250 138.150 98.210 138.605 ;
        RECT 92.320 138.105 98.210 138.150 ;
        RECT 87.865 131.965 88.285 137.015 ;
        RECT 96.630 131.965 97.050 137.015 ;
        RECT 97.710 127.025 98.210 138.105 ;
        RECT 110.125 130.540 131.985 149.320 ;
        RECT 103.900 129.990 131.985 130.540 ;
        RECT 110.125 128.920 131.985 129.990 ;
        RECT 97.710 127.010 98.665 127.025 ;
        RECT 87.870 126.510 98.665 127.010 ;
        RECT 63.755 119.725 64.145 123.095 ;
        RECT 87.870 121.960 88.290 126.510 ;
        RECT 96.630 121.960 97.050 126.510 ;
        RECT 44.895 119.350 64.145 119.725 ;
        RECT 38.245 109.855 39.530 111.910 ;
        RECT 47.970 108.660 48.870 118.430 ;
        RECT 63.755 115.930 64.145 119.350 ;
        RECT 92.250 116.160 92.670 121.210 ;
        RECT 51.835 111.360 54.335 111.700 ;
        RECT 64.125 111.370 66.625 111.710 ;
        RECT 47.920 108.105 48.920 108.660 ;
        RECT 51.835 107.800 52.735 111.360 ;
        RECT 51.785 106.875 52.780 107.800 ;
        RECT 64.125 107.175 65.025 111.370 ;
        RECT 85.625 110.385 87.210 114.270 ;
        RECT 64.075 106.250 65.075 107.175 ;
        RECT 74.615 106.020 78.035 108.380 ;
        RECT 87.885 106.330 88.375 106.880 ;
        RECT 98.115 106.000 98.665 126.510 ;
        RECT 129.345 121.845 130.955 121.870 ;
        RECT 129.345 120.285 135.250 121.845 ;
        RECT 129.345 120.260 130.955 120.285 ;
        RECT 126.765 118.495 127.185 119.145 ;
        RECT 126.760 114.115 127.180 114.765 ;
        RECT 126.540 106.330 127.180 106.880 ;
        RECT 98.115 105.450 129.030 106.000 ;
        RECT 107.220 104.280 107.795 104.830 ;
        RECT 128.480 103.950 129.030 105.450 ;
        RECT 87.920 103.400 129.030 103.950 ;
        RECT 151.760 103.135 152.760 103.900 ;
        RECT 128.675 99.590 129.605 100.140 ;
        RECT 80.585 97.560 83.555 99.105 ;
        RECT 118.360 96.880 119.570 98.825 ;
        RECT 108.185 95.255 108.605 96.005 ;
        RECT 110.765 95.255 111.185 96.005 ;
        RECT 112.225 94.655 114.120 95.030 ;
        RECT 114.495 94.655 116.390 95.030 ;
        RECT 98.875 91.320 99.295 91.905 ;
        RECT 74.615 89.460 78.030 90.575 ;
        RECT 112.690 88.740 113.160 91.790 ;
        RECT 151.815 88.260 152.705 88.285 ;
        RECT 108.735 88.100 109.235 88.125 ;
        RECT 108.735 87.735 110.660 88.100 ;
        RECT 108.735 87.710 109.235 87.735 ;
        RECT 110.280 84.565 110.660 87.735 ;
        RECT 151.810 87.360 152.710 88.260 ;
        RECT 151.815 87.335 152.705 87.360 ;
        RECT 87.440 84.185 116.860 84.565 ;
        RECT 87.440 83.515 87.820 84.185 ;
        RECT 90.020 83.515 90.400 84.185 ;
        RECT 95.180 83.515 95.560 84.185 ;
        RECT 97.760 83.515 98.140 84.185 ;
        RECT 102.920 83.515 103.300 84.185 ;
        RECT 105.500 83.515 105.880 84.185 ;
        RECT 110.660 83.515 111.040 84.185 ;
        RECT 113.240 83.510 113.620 84.185 ;
        RECT 68.150 82.640 70.495 82.665 ;
        RECT 45.055 80.285 70.500 82.640 ;
        RECT 88.710 80.635 89.130 81.685 ;
        RECT 96.450 80.635 96.870 81.685 ;
        RECT 104.190 80.635 104.610 81.685 ;
        RECT 111.930 80.635 112.350 81.685 ;
        RECT 68.150 80.260 70.495 80.285 ;
        RECT 86.150 77.150 86.850 77.160 ;
        RECT 91.310 77.150 91.690 77.160 ;
        RECT 93.890 77.150 94.270 77.160 ;
        RECT 99.050 77.150 99.430 77.160 ;
        RECT 101.630 77.150 102.010 77.160 ;
        RECT 106.790 77.150 107.170 77.160 ;
        RECT 109.370 77.150 109.750 77.160 ;
        RECT 114.530 77.150 114.910 77.160 ;
        RECT 116.490 77.150 116.860 84.185 ;
        RECT 86.150 76.780 116.860 77.150 ;
        RECT 86.150 76.110 86.530 76.780 ;
        RECT 91.310 76.110 91.690 76.780 ;
        RECT 93.890 76.110 94.270 76.780 ;
        RECT 99.050 76.110 99.430 76.780 ;
        RECT 101.630 76.110 102.010 76.780 ;
        RECT 106.790 76.110 107.170 76.780 ;
        RECT 109.370 76.110 109.750 76.780 ;
        RECT 114.530 76.110 114.910 76.780 ;
        RECT 84.840 73.230 85.260 74.280 ;
        RECT 92.580 73.230 93.000 74.280 ;
        RECT 100.320 73.230 100.740 74.280 ;
        RECT 108.060 73.230 108.480 74.280 ;
        RECT 115.800 73.230 116.220 74.280 ;
        RECT 74.615 71.055 78.035 72.090 ;
        RECT 151.760 64.430 152.760 65.165 ;
        RECT 69.765 59.435 70.890 61.390 ;
        RECT 24.335 55.870 59.430 57.795 ;
        RECT 9.465 50.075 11.565 52.125 ;
        RECT 19.090 51.320 26.875 51.690 ;
        RECT 15.540 50.630 16.590 51.050 ;
        RECT 19.090 49.740 19.460 51.320 ;
        RECT 18.420 49.360 19.470 49.740 ;
        RECT 19.090 44.580 19.460 49.360 ;
        RECT 26.495 48.450 26.875 51.320 ;
        RECT 36.965 49.325 37.340 51.220 ;
        RECT 25.820 48.070 26.875 48.450 ;
        RECT 22.945 46.760 23.995 47.180 ;
        RECT 26.495 45.870 26.875 48.070 ;
        RECT 31.050 47.520 34.100 47.990 ;
        RECT 36.965 47.055 37.340 48.950 ;
        RECT 25.825 45.490 26.875 45.870 ;
        RECT 37.565 45.595 38.315 46.015 ;
        RECT 26.495 45.110 30.410 45.490 ;
        RECT 18.420 44.200 19.470 44.580 ;
        RECT 15.540 42.890 16.590 43.310 ;
        RECT 19.090 42.000 19.460 44.200 ;
        RECT 18.420 41.620 19.470 42.000 ;
        RECT 19.090 36.840 19.460 41.620 ;
        RECT 26.495 40.710 26.875 45.110 ;
        RECT 29.985 43.780 30.410 45.110 ;
        RECT 29.960 43.280 30.435 43.780 ;
        RECT 37.565 43.015 38.315 43.435 ;
        RECT 25.825 40.330 26.875 40.710 ;
        RECT 22.945 39.020 23.995 39.440 ;
        RECT 26.495 38.130 26.875 40.330 ;
        RECT 25.825 37.750 26.875 38.130 ;
        RECT 18.420 36.460 19.470 36.840 ;
        RECT 15.540 35.150 16.590 35.570 ;
        RECT 19.090 34.260 19.460 36.460 ;
        RECT 18.420 33.880 19.470 34.260 ;
        RECT 19.090 29.100 19.460 33.880 ;
        RECT 26.495 32.970 26.875 37.750 ;
        RECT 25.825 32.590 26.875 32.970 ;
        RECT 57.505 32.795 59.430 55.870 ;
        RECT 129.460 54.995 130.730 57.045 ;
        RECT 132.440 46.490 133.440 47.315 ;
        RECT 151.760 40.410 152.760 41.175 ;
        RECT 109.100 36.505 109.490 39.875 ;
        RECT 90.240 36.130 109.490 36.505 ;
        RECT 22.945 31.280 23.995 31.700 ;
        RECT 26.495 30.390 26.875 32.590 ;
        RECT 57.480 30.820 59.455 32.795 ;
        RECT 25.825 30.010 26.875 30.390 ;
        RECT 18.420 28.720 19.470 29.100 ;
        RECT 15.540 27.410 16.590 27.830 ;
        RECT 19.090 26.520 19.460 28.720 ;
        RECT 18.420 26.140 19.470 26.520 ;
        RECT 19.090 21.680 19.460 26.140 ;
        RECT 26.495 25.230 26.875 30.010 ;
        RECT 25.825 24.850 26.875 25.230 ;
        RECT 22.945 23.540 23.995 23.960 ;
        RECT 26.495 22.650 26.875 24.850 ;
        RECT 25.825 22.270 26.875 22.650 ;
        RECT 19.090 21.360 19.470 21.680 ;
        RECT 18.420 20.980 19.470 21.360 ;
        RECT 15.540 19.670 16.590 20.090 ;
        RECT 93.315 17.855 94.215 35.210 ;
        RECT 109.100 32.710 109.490 36.130 ;
        RECT 74.530 16.955 94.215 17.855 ;
        RECT 97.180 28.140 99.680 28.480 ;
        RECT 109.470 28.150 111.970 28.490 ;
        RECT 35.840 13.265 36.840 13.860 ;
        RECT 74.530 9.090 75.430 16.955 ;
        RECT 97.180 14.025 98.080 28.140 ;
        RECT 109.470 21.505 110.370 28.150 ;
        RECT 109.420 20.605 110.420 21.505 ;
        RECT 109.470 20.595 110.370 20.605 ;
        RECT 97.130 13.125 98.130 14.025 ;
        RECT 74.480 8.190 75.480 9.090 ;
      LAYER met4 ;
        RECT 30.670 219.595 30.970 224.760 ;
        RECT 33.430 219.595 33.730 224.760 ;
        RECT 36.190 219.595 36.490 224.760 ;
        RECT 38.950 219.595 39.250 224.760 ;
        RECT 41.710 219.595 42.010 224.760 ;
        RECT 44.470 219.595 44.770 224.760 ;
        RECT 47.230 219.595 47.530 224.760 ;
        RECT 49.990 219.595 50.290 224.760 ;
        RECT 52.750 219.595 53.050 224.760 ;
        RECT 55.510 219.595 55.810 224.760 ;
        RECT 58.270 219.595 58.570 224.760 ;
        RECT 61.030 219.595 61.330 224.760 ;
        RECT 63.790 219.595 64.090 224.760 ;
        RECT 66.550 219.595 66.850 224.760 ;
        RECT 69.310 219.595 69.610 224.760 ;
        RECT 72.070 219.595 72.370 224.760 ;
        RECT 74.830 219.595 75.130 224.760 ;
        RECT 77.590 219.595 77.890 224.760 ;
        RECT 80.350 219.595 80.650 224.760 ;
        RECT 83.110 219.595 83.410 224.760 ;
        RECT 85.870 219.595 86.170 224.760 ;
        RECT 88.630 219.595 88.930 224.760 ;
        RECT 91.390 219.595 91.690 224.760 ;
        RECT 94.150 219.595 94.450 224.760 ;
        RECT 4.000 216.410 95.080 219.595 ;
        RECT 85.690 152.800 87.500 152.810 ;
        RECT 80.155 150.800 157.000 152.800 ;
        RECT 80.155 149.315 99.300 150.800 ;
        RECT 80.155 138.890 83.640 149.315 ;
        RECT 86.110 148.275 99.300 149.315 ;
        RECT 87.910 132.485 88.240 136.995 ;
        RECT 96.675 132.485 97.005 136.995 ;
        RECT 87.910 131.985 100.180 132.485 ;
        RECT 92.295 121.015 92.625 121.190 ;
        RECT 99.680 121.015 100.180 131.985 ;
        RECT 110.520 129.315 130.130 148.925 ;
        RECT 92.295 120.515 100.180 121.015 ;
        RECT 92.295 116.180 92.625 120.515 ;
        RECT 85.670 114.245 87.165 114.250 ;
        RECT 38.290 111.885 39.485 111.890 ;
        RECT 4.000 109.880 39.485 111.885 ;
        RECT 80.630 110.410 87.165 114.245 ;
        RECT 80.630 110.405 83.445 110.410 ;
        RECT 85.670 110.405 87.165 110.410 ;
        RECT 38.290 109.875 39.485 109.880 ;
        RECT 51.830 106.870 52.735 107.805 ;
        RECT 45.080 82.640 47.445 82.645 ;
        RECT 4.000 80.285 47.445 82.640 ;
        RECT 45.080 80.280 47.445 80.285 ;
        RECT 24.360 57.795 26.295 57.800 ;
        RECT 4.000 55.870 26.295 57.795 ;
        RECT 24.360 55.865 26.295 55.870 ;
        RECT 19.215 52.980 37.330 53.360 ;
        RECT 19.215 52.420 19.600 52.980 ;
        RECT 9.510 52.100 11.520 52.105 ;
        RECT 4.000 50.100 11.520 52.100 ;
        RECT 9.510 50.095 11.520 50.100 ;
        RECT 15.560 52.040 23.345 52.420 ;
        RECT 15.560 51.005 15.940 52.040 ;
        RECT 15.560 50.675 16.570 51.005 ;
        RECT 15.560 43.265 15.940 50.675 ;
        RECT 22.965 47.135 23.345 52.040 ;
        RECT 31.070 47.565 34.100 47.945 ;
        RECT 22.965 46.805 23.975 47.135 ;
        RECT 15.560 42.935 16.570 43.265 ;
        RECT 15.560 35.525 15.940 42.935 ;
        RECT 22.965 39.395 23.345 46.805 ;
        RECT 33.720 44.665 34.100 47.565 ;
        RECT 36.965 46.915 37.330 52.980 ;
        RECT 36.060 45.640 38.295 45.970 ;
        RECT 36.060 44.665 36.440 45.640 ;
        RECT 33.720 44.335 36.440 44.665 ;
        RECT 36.060 43.390 36.440 44.335 ;
        RECT 36.060 43.060 38.295 43.390 ;
        RECT 22.965 39.065 23.975 39.395 ;
        RECT 15.560 35.195 16.570 35.525 ;
        RECT 15.560 27.785 15.940 35.195 ;
        RECT 22.965 31.655 23.345 39.065 ;
        RECT 22.965 31.325 23.975 31.655 ;
        RECT 15.560 27.455 16.570 27.785 ;
        RECT 15.560 20.045 15.940 27.455 ;
        RECT 22.965 23.915 23.345 31.325 ;
        RECT 22.965 23.585 23.975 23.915 ;
        RECT 15.560 19.715 16.570 20.045 ;
        RECT 51.835 14.025 52.735 106.870 ;
        RECT 64.120 106.245 65.030 107.180 ;
        RECT 64.125 21.505 65.025 106.245 ;
        RECT 74.660 106.040 77.990 108.360 ;
        RECT 74.665 90.555 77.985 106.040 ;
        RECT 80.635 99.085 83.445 110.405 ;
        RECT 99.680 106.860 100.180 120.515 ;
        RECT 126.810 118.515 127.140 129.315 ;
        RECT 131.485 128.980 131.965 149.260 ;
        RECT 133.655 121.845 135.225 121.850 ;
        RECT 133.655 120.285 157.000 121.845 ;
        RECT 133.655 120.280 135.225 120.285 ;
        RECT 126.805 106.860 127.135 114.745 ;
        RECT 87.965 106.350 130.370 106.860 ;
        RECT 129.860 106.160 130.370 106.350 ;
        RECT 129.860 105.260 152.710 106.160 ;
        RECT 129.860 104.810 130.370 105.260 ;
        RECT 107.345 104.300 130.370 104.810 ;
        RECT 151.810 103.880 152.710 105.260 ;
        RECT 151.805 103.155 152.715 103.880 ;
        RECT 128.720 100.115 129.560 100.120 ;
        RECT 98.920 99.615 129.560 100.115 ;
        RECT 80.630 97.580 83.510 99.085 ;
        RECT 98.920 91.340 99.250 99.615 ;
        RECT 128.720 99.610 129.560 99.615 ;
        RECT 118.405 98.800 119.525 98.805 ;
        RECT 118.405 96.905 157.000 98.800 ;
        RECT 118.405 96.900 119.525 96.905 ;
        RECT 108.230 94.130 108.560 95.985 ;
        RECT 110.810 94.130 111.140 95.985 ;
        RECT 112.085 94.655 118.530 95.020 ;
        RECT 108.230 93.750 111.140 94.130 ;
        RECT 109.505 91.790 109.835 93.750 ;
        RECT 109.505 91.410 113.115 91.790 ;
        RECT 74.660 89.480 77.985 90.555 ;
        RECT 74.665 82.640 77.985 89.480 ;
        RECT 112.735 88.760 113.115 91.410 ;
        RECT 68.145 80.285 77.985 82.640 ;
        RECT 88.755 81.035 89.085 81.665 ;
        RECT 96.495 81.035 96.825 81.665 ;
        RECT 104.235 81.035 104.565 81.665 ;
        RECT 111.975 81.035 112.305 81.665 ;
        RECT 88.755 80.655 117.590 81.035 ;
        RECT 74.665 72.070 77.985 80.285 ;
        RECT 117.210 77.290 117.590 80.655 ;
        RECT 118.150 77.290 118.530 94.655 ;
        RECT 117.210 76.905 118.530 77.290 ;
        RECT 84.885 73.630 85.215 74.260 ;
        RECT 92.625 73.630 92.955 74.260 ;
        RECT 100.365 73.630 100.695 74.260 ;
        RECT 108.105 73.630 108.435 74.260 ;
        RECT 115.845 73.630 116.175 74.260 ;
        RECT 117.210 73.630 117.590 76.905 ;
        RECT 84.885 73.250 117.590 73.630 ;
        RECT 74.660 71.075 77.990 72.070 ;
        RECT 151.810 65.145 152.710 88.260 ;
        RECT 151.805 64.450 152.715 65.145 ;
        RECT 69.810 61.365 70.845 61.370 ;
        RECT 69.810 59.460 139.665 61.365 ;
        RECT 69.810 59.455 70.845 59.460 ;
        RECT 129.505 57.020 130.685 57.025 ;
        RECT 137.760 57.020 139.665 59.460 ;
        RECT 129.505 55.020 157.000 57.020 ;
        RECT 129.505 55.015 130.685 55.020 ;
        RECT 132.485 46.510 133.395 47.295 ;
        RECT 109.465 21.505 110.375 21.510 ;
        RECT 64.125 20.605 114.070 21.505 ;
        RECT 109.465 20.600 110.375 20.605 ;
        RECT 97.175 14.025 98.085 14.030 ;
        RECT 35.885 13.285 36.795 13.840 ;
        RECT 35.890 8.415 36.790 13.285 ;
        RECT 51.835 13.125 98.085 14.025 ;
        RECT 35.890 7.515 56.110 8.415 ;
        RECT 74.525 8.185 75.435 9.095 ;
        RECT 55.210 1.690 56.110 7.515 ;
        RECT 55.205 1.000 56.110 1.690 ;
        RECT 74.530 1.000 75.430 8.185 ;
        RECT 93.850 1.000 94.750 13.125 ;
        RECT 97.175 13.120 98.085 13.125 ;
        RECT 113.170 1.000 114.070 20.605 ;
        RECT 132.490 1.000 133.390 46.510 ;
        RECT 151.805 40.430 152.715 41.155 ;
        RECT 151.810 1.000 152.710 40.430 ;
        RECT 55.205 0.995 55.210 1.000 ;
  END
END tt_um_DalinEM_diff_amp
END LIBRARY

