magic
tech sky130A
magscale 1 2
timestamp 1738877391
<< nwell >>
rect -437 1479 275 2117
rect 853 1479 1565 2117
rect 2143 1479 2855 2117
rect 3404 1459 4739 2338
<< pwell >>
rect -928 587 4746 1434
<< pmoslvt >>
rect -241 1698 79 1898
rect 1049 1698 1369 1898
rect 2339 1698 2659 1898
rect 3629 1698 3949 1898
rect 4265 1698 4465 1898
<< nmoslvt >>
rect -637 911 -437 1111
rect -379 911 -179 1111
rect -121 911 79 1111
rect 137 911 337 1111
rect 395 911 595 1111
rect 653 911 853 1111
rect 911 911 1111 1111
rect 1169 911 1369 1111
rect 1427 911 1627 1111
rect 1685 911 1885 1111
rect 1943 911 2143 1111
rect 2201 911 2401 1111
rect 2459 911 2659 1111
rect 2717 911 2917 1111
rect 2975 911 3175 1111
rect 3233 911 3433 1111
rect 3491 911 3691 1111
rect 3749 911 3949 1111
rect 4007 911 4207 1111
rect 4265 911 4465 1111
<< ndiff >>
rect -695 1099 -637 1111
rect -695 923 -683 1099
rect -649 923 -637 1099
rect -695 911 -637 923
rect -437 1099 -379 1111
rect -437 923 -425 1099
rect -391 923 -379 1099
rect -437 911 -379 923
rect -179 1099 -121 1111
rect -179 923 -167 1099
rect -133 923 -121 1099
rect -179 911 -121 923
rect 79 1099 137 1111
rect 79 923 91 1099
rect 125 923 137 1099
rect 79 911 137 923
rect 337 1099 395 1111
rect 337 923 349 1099
rect 383 923 395 1099
rect 337 911 395 923
rect 595 1099 653 1111
rect 595 923 607 1099
rect 641 923 653 1099
rect 595 911 653 923
rect 853 1099 911 1111
rect 853 923 865 1099
rect 899 923 911 1099
rect 853 911 911 923
rect 1111 1099 1169 1111
rect 1111 923 1123 1099
rect 1157 923 1169 1099
rect 1111 911 1169 923
rect 1369 1099 1427 1111
rect 1369 923 1381 1099
rect 1415 923 1427 1099
rect 1369 911 1427 923
rect 1627 1099 1685 1111
rect 1627 923 1639 1099
rect 1673 923 1685 1099
rect 1627 911 1685 923
rect 1885 1099 1943 1111
rect 1885 923 1897 1099
rect 1931 923 1943 1099
rect 1885 911 1943 923
rect 2143 1099 2201 1111
rect 2143 923 2155 1099
rect 2189 923 2201 1099
rect 2143 911 2201 923
rect 2401 1099 2459 1111
rect 2401 923 2413 1099
rect 2447 923 2459 1099
rect 2401 911 2459 923
rect 2659 1099 2717 1111
rect 2659 923 2671 1099
rect 2705 923 2717 1099
rect 2659 911 2717 923
rect 2917 1099 2975 1111
rect 2917 923 2929 1099
rect 2963 923 2975 1099
rect 2917 911 2975 923
rect 3175 1099 3233 1111
rect 3175 923 3187 1099
rect 3221 923 3233 1099
rect 3175 911 3233 923
rect 3433 1099 3491 1111
rect 3433 923 3445 1099
rect 3479 923 3491 1099
rect 3433 911 3491 923
rect 3691 1099 3749 1111
rect 3691 923 3703 1099
rect 3737 923 3749 1099
rect 3691 911 3749 923
rect 3949 1099 4007 1111
rect 3949 923 3961 1099
rect 3995 923 4007 1099
rect 3949 911 4007 923
rect 4207 1099 4265 1111
rect 4207 923 4219 1099
rect 4253 923 4265 1099
rect 4207 911 4265 923
rect 4465 1099 4523 1111
rect 4465 923 4477 1099
rect 4511 923 4523 1099
rect 4465 911 4523 923
<< pdiff >>
rect -299 1886 -241 1898
rect -299 1710 -287 1886
rect -253 1710 -241 1886
rect -299 1698 -241 1710
rect 79 1886 137 1898
rect 79 1710 91 1886
rect 125 1710 137 1886
rect 79 1698 137 1710
rect 991 1886 1049 1898
rect 991 1710 1003 1886
rect 1037 1710 1049 1886
rect 991 1698 1049 1710
rect 1369 1886 1427 1898
rect 1369 1710 1381 1886
rect 1415 1710 1427 1886
rect 1369 1698 1427 1710
rect 2281 1886 2339 1898
rect 2281 1710 2293 1886
rect 2327 1710 2339 1886
rect 2281 1698 2339 1710
rect 2659 1886 2717 1898
rect 2659 1710 2671 1886
rect 2705 1710 2717 1886
rect 2659 1698 2717 1710
rect 3571 1886 3629 1898
rect 3571 1710 3583 1886
rect 3617 1710 3629 1886
rect 3571 1698 3629 1710
rect 3949 1886 4007 1898
rect 3949 1710 3961 1886
rect 3995 1710 4007 1886
rect 3949 1698 4007 1710
rect 4207 1886 4265 1898
rect 4207 1710 4219 1886
rect 4253 1710 4265 1886
rect 4207 1698 4265 1710
rect 4465 1886 4523 1898
rect 4465 1710 4477 1886
rect 4511 1710 4523 1886
rect 4465 1698 4523 1710
<< ndiffc >>
rect -683 923 -649 1099
rect -425 923 -391 1099
rect -167 923 -133 1099
rect 91 923 125 1099
rect 349 923 383 1099
rect 607 923 641 1099
rect 865 923 899 1099
rect 1123 923 1157 1099
rect 1381 923 1415 1099
rect 1639 923 1673 1099
rect 1897 923 1931 1099
rect 2155 923 2189 1099
rect 2413 923 2447 1099
rect 2671 923 2705 1099
rect 2929 923 2963 1099
rect 3187 923 3221 1099
rect 3445 923 3479 1099
rect 3703 923 3737 1099
rect 3961 923 3995 1099
rect 4219 923 4253 1099
rect 4477 923 4511 1099
<< pdiffc >>
rect -287 1710 -253 1886
rect 91 1710 125 1886
rect 1003 1710 1037 1886
rect 1381 1710 1415 1886
rect 2293 1710 2327 1886
rect 2671 1710 2705 1886
rect 3583 1710 3617 1886
rect 3961 1710 3995 1886
rect 4219 1710 4253 1886
rect 4477 1710 4511 1886
<< psubdiff >>
rect -850 1333 -790 1367
rect 4618 1333 4678 1367
rect -850 1307 -816 1333
rect 4644 1307 4678 1333
rect -850 699 -816 725
rect 4644 699 4678 725
rect -850 665 -790 699
rect 4618 665 4678 699
<< nsubdiff >>
rect 3472 2260 3532 2294
rect 4598 2260 4658 2294
rect 3472 2206 3506 2260
rect -401 2047 -305 2081
rect 143 2047 239 2081
rect -401 1985 -367 2047
rect 205 1985 239 2047
rect -401 1549 -367 1611
rect 205 1549 239 1611
rect -401 1515 -305 1549
rect 143 1515 239 1549
rect 889 2047 985 2081
rect 1433 2047 1529 2081
rect 889 1985 923 2047
rect 1495 1985 1529 2047
rect 889 1549 923 1611
rect 1495 1549 1529 1611
rect 889 1515 985 1549
rect 1433 1515 1529 1549
rect 2179 2047 2275 2081
rect 2723 2047 2819 2081
rect 2179 1985 2213 2047
rect 2785 1985 2819 2047
rect 2179 1549 2213 1611
rect 2785 1549 2819 1611
rect 2179 1515 2275 1549
rect 2723 1515 2819 1549
rect 4624 2206 4658 2260
rect 3472 1556 3506 1582
rect 4624 1556 4658 1582
rect 3472 1522 3532 1556
rect 4598 1522 4658 1556
<< psubdiffcont >>
rect -790 1333 4618 1367
rect -850 725 -816 1307
rect 4644 725 4678 1307
rect -790 665 4618 699
<< nsubdiffcont >>
rect 3532 2260 4598 2294
rect -305 2047 143 2081
rect -401 1611 -367 1985
rect 205 1611 239 1985
rect -305 1515 143 1549
rect 985 2047 1433 2081
rect 889 1611 923 1985
rect 1495 1611 1529 1985
rect 985 1515 1433 1549
rect 2275 2047 2723 2081
rect 2179 1611 2213 1985
rect 2785 1611 2819 1985
rect 2275 1515 2723 1549
rect 3472 1582 3506 2206
rect 4624 1582 4658 2206
rect 3532 1522 4598 1556
<< poly >>
rect -241 1979 79 1995
rect -241 1945 -225 1979
rect 63 1945 79 1979
rect -241 1898 79 1945
rect -241 1651 79 1698
rect -241 1617 -225 1651
rect 63 1617 79 1651
rect -241 1601 79 1617
rect 1049 1979 1369 1995
rect 1049 1945 1065 1979
rect 1353 1945 1369 1979
rect 1049 1898 1369 1945
rect 1049 1651 1369 1698
rect 1049 1617 1065 1651
rect 1353 1617 1369 1651
rect 1049 1601 1369 1617
rect 2339 1979 2659 1995
rect 2339 1945 2355 1979
rect 2643 1945 2659 1979
rect 2339 1898 2659 1945
rect 2339 1651 2659 1698
rect 2339 1617 2355 1651
rect 2643 1617 2659 1651
rect 2339 1601 2659 1617
rect 3629 1979 3949 1995
rect 3629 1945 3645 1979
rect 3933 1945 3949 1979
rect 3629 1898 3949 1945
rect 4265 1979 4465 1995
rect 4265 1945 4281 1979
rect 4449 1945 4465 1979
rect 4265 1898 4465 1945
rect 3629 1651 3949 1698
rect 3629 1617 3645 1651
rect 3933 1617 3949 1651
rect 3629 1601 3949 1617
rect 4265 1651 4465 1698
rect 4265 1617 4281 1651
rect 4449 1617 4465 1651
rect 4265 1601 4465 1617
rect -637 1183 -437 1199
rect -637 1149 -621 1183
rect -453 1149 -437 1183
rect -637 1111 -437 1149
rect -379 1183 -179 1199
rect -379 1149 -363 1183
rect -195 1149 -179 1183
rect -379 1111 -179 1149
rect -121 1183 79 1199
rect -121 1149 -105 1183
rect 63 1149 79 1183
rect -121 1111 79 1149
rect 137 1183 337 1199
rect 137 1149 153 1183
rect 321 1149 337 1183
rect 137 1111 337 1149
rect 395 1183 595 1199
rect 395 1149 411 1183
rect 579 1149 595 1183
rect 395 1111 595 1149
rect 653 1183 853 1199
rect 653 1149 669 1183
rect 837 1149 853 1183
rect 653 1111 853 1149
rect 911 1183 1111 1199
rect 911 1149 927 1183
rect 1095 1149 1111 1183
rect 911 1111 1111 1149
rect 1169 1183 1369 1199
rect 1169 1149 1185 1183
rect 1353 1149 1369 1183
rect 1169 1111 1369 1149
rect 1427 1183 1627 1199
rect 1427 1149 1443 1183
rect 1611 1149 1627 1183
rect 1427 1111 1627 1149
rect 1685 1183 1885 1199
rect 1685 1149 1701 1183
rect 1869 1149 1885 1183
rect 1685 1111 1885 1149
rect 1943 1183 2143 1199
rect 1943 1149 1959 1183
rect 2127 1149 2143 1183
rect 1943 1111 2143 1149
rect 2201 1183 2401 1199
rect 2201 1149 2217 1183
rect 2385 1149 2401 1183
rect 2201 1111 2401 1149
rect 2459 1183 2659 1199
rect 2459 1149 2475 1183
rect 2643 1149 2659 1183
rect 2459 1111 2659 1149
rect 2717 1183 2917 1199
rect 2717 1149 2733 1183
rect 2901 1149 2917 1183
rect 2717 1111 2917 1149
rect 2975 1183 3175 1199
rect 2975 1149 2991 1183
rect 3159 1149 3175 1183
rect 2975 1111 3175 1149
rect 3233 1183 3433 1199
rect 3233 1149 3249 1183
rect 3417 1149 3433 1183
rect 3233 1111 3433 1149
rect 3491 1183 3691 1199
rect 3491 1149 3507 1183
rect 3675 1149 3691 1183
rect 3491 1111 3691 1149
rect 3749 1183 3949 1199
rect 3749 1149 3765 1183
rect 3933 1149 3949 1183
rect 3749 1111 3949 1149
rect 4007 1183 4207 1199
rect 4007 1149 4023 1183
rect 4191 1149 4207 1183
rect 4007 1111 4207 1149
rect 4265 1183 4465 1199
rect 4265 1149 4281 1183
rect 4449 1149 4465 1183
rect 4265 1111 4465 1149
rect -637 873 -437 911
rect -637 839 -621 873
rect -453 839 -437 873
rect -637 823 -437 839
rect -379 873 -179 911
rect -379 839 -363 873
rect -195 839 -179 873
rect -379 823 -179 839
rect -121 873 79 911
rect -121 839 -105 873
rect 63 839 79 873
rect -121 823 79 839
rect 137 873 337 911
rect 137 839 153 873
rect 321 839 337 873
rect 137 823 337 839
rect 395 873 595 911
rect 395 839 411 873
rect 579 839 595 873
rect 395 823 595 839
rect 653 873 853 911
rect 653 839 669 873
rect 837 839 853 873
rect 653 823 853 839
rect 911 873 1111 911
rect 911 839 927 873
rect 1095 839 1111 873
rect 911 823 1111 839
rect 1169 873 1369 911
rect 1169 839 1185 873
rect 1353 839 1369 873
rect 1169 823 1369 839
rect 1427 873 1627 911
rect 1427 839 1443 873
rect 1611 839 1627 873
rect 1427 823 1627 839
rect 1685 873 1885 911
rect 1685 839 1701 873
rect 1869 839 1885 873
rect 1685 823 1885 839
rect 1943 873 2143 911
rect 1943 839 1959 873
rect 2127 839 2143 873
rect 1943 823 2143 839
rect 2201 873 2401 911
rect 2201 839 2217 873
rect 2385 839 2401 873
rect 2201 823 2401 839
rect 2459 873 2659 911
rect 2459 839 2475 873
rect 2643 839 2659 873
rect 2459 823 2659 839
rect 2717 873 2917 911
rect 2717 839 2733 873
rect 2901 839 2917 873
rect 2717 823 2917 839
rect 2975 873 3175 911
rect 2975 839 2991 873
rect 3159 839 3175 873
rect 2975 823 3175 839
rect 3233 873 3433 911
rect 3233 839 3249 873
rect 3417 839 3433 873
rect 3233 823 3433 839
rect 3491 873 3691 911
rect 3491 839 3507 873
rect 3675 839 3691 873
rect 3491 823 3691 839
rect 3749 873 3949 911
rect 3749 839 3765 873
rect 3933 839 3949 873
rect 3749 823 3949 839
rect 4007 873 4207 911
rect 4007 839 4023 873
rect 4191 839 4207 873
rect 4007 823 4207 839
rect 4265 873 4465 911
rect 4265 839 4281 873
rect 4449 839 4465 873
rect 4265 823 4465 839
<< polycont >>
rect -225 1945 63 1979
rect -225 1617 63 1651
rect 1065 1945 1353 1979
rect 1065 1617 1353 1651
rect 2355 1945 2643 1979
rect 2355 1617 2643 1651
rect 3645 1945 3933 1979
rect 4281 1945 4449 1979
rect 3645 1617 3933 1651
rect 4281 1617 4449 1651
rect -621 1149 -453 1183
rect -363 1149 -195 1183
rect -105 1149 63 1183
rect 153 1149 321 1183
rect 411 1149 579 1183
rect 669 1149 837 1183
rect 927 1149 1095 1183
rect 1185 1149 1353 1183
rect 1443 1149 1611 1183
rect 1701 1149 1869 1183
rect 1959 1149 2127 1183
rect 2217 1149 2385 1183
rect 2475 1149 2643 1183
rect 2733 1149 2901 1183
rect 2991 1149 3159 1183
rect 3249 1149 3417 1183
rect 3507 1149 3675 1183
rect 3765 1149 3933 1183
rect 4023 1149 4191 1183
rect 4281 1149 4449 1183
rect -621 839 -453 873
rect -363 839 -195 873
rect -105 839 63 873
rect 153 839 321 873
rect 411 839 579 873
rect 669 839 837 873
rect 927 839 1095 873
rect 1185 839 1353 873
rect 1443 839 1611 873
rect 1701 839 1869 873
rect 1959 839 2127 873
rect 2217 839 2385 873
rect 2475 839 2643 873
rect 2733 839 2901 873
rect 2991 839 3159 873
rect 3249 839 3417 873
rect 3507 839 3675 873
rect 3765 839 3933 873
rect 4023 839 4191 873
rect 4281 839 4449 873
<< locali >>
rect -423 2296 4741 2352
rect -423 2157 -374 2296
rect -423 2081 3472 2157
rect -423 2047 -305 2081
rect 143 2047 985 2081
rect 1433 2047 2275 2081
rect 2723 2047 3472 2081
rect -423 2027 3472 2047
rect -423 1985 -329 2027
rect -423 1611 -401 1985
rect -367 1611 -329 1985
rect 177 1985 278 2027
rect -241 1945 -225 1979
rect 63 1945 79 1979
rect -287 1886 -253 1902
rect -287 1694 -253 1710
rect 91 1886 125 1902
rect 91 1694 125 1710
rect -241 1617 -225 1651
rect 63 1617 79 1651
rect -423 1576 -329 1611
rect 177 1611 205 1985
rect 239 1611 278 1985
rect 177 1576 278 1611
rect -423 1549 278 1576
rect -423 1515 -305 1549
rect 143 1515 278 1549
rect -423 1479 278 1515
rect 852 1985 968 2027
rect 852 1611 889 1985
rect 923 1611 968 1985
rect 1465 1985 1572 2027
rect 1049 1945 1065 1979
rect 1353 1945 1369 1979
rect 1003 1886 1037 1902
rect 1003 1694 1037 1710
rect 1381 1886 1415 1902
rect 1381 1694 1415 1710
rect 1049 1617 1065 1651
rect 1353 1617 1369 1651
rect 852 1573 968 1611
rect 1465 1611 1495 1985
rect 1529 1611 1572 1985
rect 1465 1573 1572 1611
rect 852 1549 1572 1573
rect 852 1515 985 1549
rect 1433 1515 1572 1549
rect 852 1476 1572 1515
rect 2165 1985 2258 2027
rect 2165 1611 2179 1985
rect 2213 1611 2258 1985
rect 2758 1985 2865 2027
rect 3364 2023 3472 2027
rect 2339 1945 2355 1979
rect 2643 1945 2659 1979
rect 2293 1886 2327 1902
rect 2293 1694 2327 1710
rect 2671 1886 2705 1902
rect 2671 1694 2705 1710
rect 2339 1617 2355 1651
rect 2643 1617 2659 1651
rect 2165 1577 2258 1611
rect 2758 1611 2785 1985
rect 2819 1611 2865 1985
rect 2758 1577 2865 1611
rect 2165 1549 2865 1577
rect 2165 1515 2275 1549
rect 2723 1515 2865 1549
rect 2165 1480 2865 1515
rect 3404 1582 3472 2023
rect 3506 2023 4624 2157
rect 3506 1582 3530 2023
rect 3629 1945 3645 1979
rect 3933 1945 3949 1979
rect 4265 1945 4281 1979
rect 4449 1945 4465 1979
rect 3583 1886 3617 1902
rect 3583 1694 3617 1710
rect 3961 1886 3995 1902
rect 3961 1694 3995 1710
rect 4219 1886 4253 1902
rect 4219 1694 4253 1710
rect 4477 1886 4511 1902
rect 4477 1694 4511 1710
rect 3629 1617 3645 1651
rect 3933 1617 3949 1651
rect 4265 1617 4281 1651
rect 4449 1617 4465 1651
rect 3404 1572 3530 1582
rect 4598 1582 4624 2023
rect 4658 1582 4741 2296
rect 4598 1572 4741 1582
rect 3404 1563 4741 1572
rect 3404 1556 4740 1563
rect 3404 1522 3532 1556
rect 4598 1522 4740 1556
rect 3404 1459 4740 1522
rect -897 1367 4725 1425
rect -897 1333 -790 1367
rect 4618 1333 4725 1367
rect -897 1307 4725 1333
rect -897 725 -850 1307
rect -816 1286 4644 1307
rect -816 791 -774 1286
rect -637 1149 -621 1183
rect -453 1149 -437 1183
rect -379 1149 -363 1183
rect -195 1149 -179 1183
rect -121 1149 -105 1183
rect 63 1149 79 1183
rect 137 1149 153 1183
rect 321 1149 337 1183
rect 395 1149 411 1183
rect 579 1149 595 1183
rect 653 1149 669 1183
rect 837 1149 853 1183
rect 911 1149 927 1183
rect 1095 1149 1111 1183
rect 1169 1149 1185 1183
rect 1353 1149 1369 1183
rect 1427 1149 1443 1183
rect 1611 1149 1627 1183
rect 1685 1149 1701 1183
rect 1869 1149 1885 1183
rect 1943 1149 1959 1183
rect 2127 1149 2143 1183
rect 2201 1149 2217 1183
rect 2385 1149 2401 1183
rect 2459 1149 2475 1183
rect 2643 1149 2659 1183
rect 2717 1149 2733 1183
rect 2901 1149 2917 1183
rect 2975 1149 2991 1183
rect 3159 1149 3175 1183
rect 3233 1149 3249 1183
rect 3417 1149 3433 1183
rect 3491 1149 3507 1183
rect 3675 1149 3691 1183
rect 3749 1149 3765 1183
rect 3933 1149 3949 1183
rect 4007 1149 4023 1183
rect 4191 1149 4207 1183
rect 4265 1149 4281 1183
rect 4449 1149 4465 1183
rect -683 1099 -649 1115
rect -683 907 -649 923
rect -425 1099 -391 1115
rect -425 907 -391 923
rect -167 1099 -133 1115
rect -167 907 -133 923
rect 91 1099 125 1115
rect 91 907 125 923
rect 349 1099 383 1115
rect 349 907 383 923
rect 607 1099 641 1115
rect 607 907 641 923
rect 865 1099 899 1115
rect 865 907 899 923
rect 1123 1099 1157 1115
rect 1123 907 1157 923
rect 1381 1099 1415 1115
rect 1381 907 1415 923
rect 1639 1099 1673 1115
rect 1639 907 1673 923
rect 1897 1099 1931 1115
rect 1897 907 1931 923
rect 2155 1099 2189 1115
rect 2155 907 2189 923
rect 2413 1099 2447 1115
rect 2413 907 2447 923
rect 2671 1099 2705 1115
rect 2671 907 2705 923
rect 2929 1099 2963 1115
rect 2929 907 2963 923
rect 3187 1099 3221 1115
rect 3187 907 3221 923
rect 3445 1099 3479 1115
rect 3445 907 3479 923
rect 3703 1099 3737 1115
rect 3703 907 3737 923
rect 3961 1099 3995 1115
rect 3961 907 3995 923
rect 4219 1099 4253 1115
rect 4219 907 4253 923
rect 4477 1099 4511 1115
rect 4477 907 4511 923
rect -637 839 -621 873
rect -453 839 -437 873
rect -379 839 -363 873
rect -195 839 -179 873
rect -121 839 -105 873
rect 63 839 79 873
rect 137 839 153 873
rect 321 839 337 873
rect 395 839 411 873
rect 579 839 595 873
rect 653 839 669 873
rect 837 839 853 873
rect 911 839 927 873
rect 1095 839 1111 873
rect 1169 839 1185 873
rect 1353 839 1369 873
rect 1427 839 1443 873
rect 1611 839 1627 873
rect 1685 839 1701 873
rect 1869 839 1885 873
rect 1943 839 1959 873
rect 2127 839 2143 873
rect 2201 839 2217 873
rect 2385 839 2401 873
rect 2459 839 2475 873
rect 2643 839 2659 873
rect 2717 839 2733 873
rect 2901 839 2917 873
rect 2975 839 2991 873
rect 3159 839 3175 873
rect 3233 839 3249 873
rect 3417 839 3433 873
rect 3491 839 3507 873
rect 3675 839 3691 873
rect 3749 839 3765 873
rect 3933 839 3949 873
rect 4007 839 4023 873
rect 4191 839 4207 873
rect 4265 839 4281 873
rect 4449 839 4465 873
rect 4602 791 4644 1286
rect -816 754 4644 791
rect -816 725 -804 754
rect -897 563 -804 725
rect 4603 725 4644 754
rect 4678 725 4725 1307
rect 4603 699 4725 725
rect 4618 665 4725 699
rect 4603 563 4725 665
rect -897 535 4725 563
<< viali >>
rect -374 2294 4658 2296
rect -374 2260 3532 2294
rect 3532 2260 4598 2294
rect 4598 2260 4658 2294
rect -374 2206 4658 2260
rect -374 2157 3472 2206
rect 3472 2157 3506 2206
rect 3506 2157 4624 2206
rect 4624 2157 4658 2206
rect -225 1945 63 1979
rect -287 1710 -253 1886
rect 91 1710 125 1886
rect -225 1617 63 1651
rect 1065 1945 1353 1979
rect 1003 1710 1037 1886
rect 1381 1710 1415 1886
rect 1065 1617 1353 1651
rect 2355 1945 2643 1979
rect 2293 1710 2327 1886
rect 2671 1710 2705 1886
rect 2355 1617 2643 1651
rect 3645 1945 3933 1979
rect 4281 1945 4449 1979
rect 3583 1710 3617 1886
rect 3961 1710 3995 1886
rect 4219 1710 4253 1886
rect 4477 1710 4511 1886
rect 3645 1617 3933 1651
rect 4281 1617 4449 1651
rect -621 1149 -453 1183
rect -363 1149 -195 1183
rect -105 1149 63 1183
rect 153 1149 321 1183
rect 411 1149 579 1183
rect 669 1149 837 1183
rect 927 1149 1095 1183
rect 1185 1149 1353 1183
rect 1443 1149 1611 1183
rect 1701 1149 1869 1183
rect 1959 1149 2127 1183
rect 2217 1149 2385 1183
rect 2475 1149 2643 1183
rect 2733 1149 2901 1183
rect 2991 1149 3159 1183
rect 3249 1149 3417 1183
rect 3507 1149 3675 1183
rect 3765 1149 3933 1183
rect 4023 1149 4191 1183
rect 4281 1149 4449 1183
rect -683 923 -649 1099
rect -425 923 -391 1099
rect -167 923 -133 1099
rect 91 923 125 1099
rect 349 923 383 1099
rect 607 923 641 1099
rect 865 923 899 1099
rect 1123 923 1157 1099
rect 1381 923 1415 1099
rect 1639 923 1673 1099
rect 1897 923 1931 1099
rect 2155 923 2189 1099
rect 2413 923 2447 1099
rect 2671 923 2705 1099
rect 2929 923 2963 1099
rect 3187 923 3221 1099
rect 3445 923 3479 1099
rect 3703 923 3737 1099
rect 3961 923 3995 1099
rect 4219 923 4253 1099
rect 4477 923 4511 1099
rect -621 839 -453 873
rect -363 839 -195 873
rect -105 839 63 873
rect 153 839 321 873
rect 411 839 579 873
rect 669 839 837 873
rect 927 839 1095 873
rect 1185 839 1353 873
rect 1443 839 1611 873
rect 1701 839 1869 873
rect 1959 839 2127 873
rect 2217 839 2385 873
rect 2475 839 2643 873
rect 2733 839 2901 873
rect 2991 839 3159 873
rect 3249 839 3417 873
rect 3507 839 3675 873
rect 3765 839 3933 873
rect 4023 839 4191 873
rect 4281 839 4449 873
rect -804 699 4603 754
rect -804 665 -790 699
rect -790 665 4603 699
rect -804 563 4603 665
<< metal1 >>
rect -386 2296 4670 2302
rect -386 2157 -374 2296
rect 4658 2157 4670 2296
rect -386 2151 4670 2157
rect -237 1979 75 1985
rect -237 1945 -225 1979
rect 63 1945 75 1979
rect -237 1939 75 1945
rect 1053 1979 1365 1985
rect 1053 1945 1065 1979
rect 1353 1945 1365 1979
rect 1053 1939 1365 1945
rect 2343 1979 2655 1985
rect 2343 1945 2355 1979
rect 2643 1945 2655 1979
rect 2343 1939 2655 1945
rect 3633 1979 3945 1985
rect 3633 1945 3645 1979
rect 3933 1945 3945 1979
rect 3633 1939 3945 1945
rect 4269 1979 4461 1985
rect 4269 1945 4281 1979
rect 4449 1945 4461 1979
rect 4269 1939 4461 1945
rect -293 1886 -247 1898
rect -306 1826 -296 1886
rect -244 1826 -234 1886
rect -293 1710 -287 1826
rect -253 1710 -247 1826
rect -293 1698 -247 1710
rect -164 1657 11 1939
rect 85 1886 131 1898
rect 997 1886 1043 1898
rect 85 1770 91 1886
rect 125 1770 131 1886
rect 984 1816 994 1886
rect 1046 1816 1056 1886
rect 72 1710 82 1770
rect 134 1710 144 1770
rect 997 1710 1003 1816
rect 1037 1710 1043 1816
rect 85 1698 131 1710
rect 997 1698 1043 1710
rect 1132 1657 1307 1939
rect 1375 1886 1421 1898
rect 2287 1886 2333 1898
rect 1375 1780 1381 1886
rect 1415 1780 1421 1886
rect 2274 1816 2284 1886
rect 2336 1816 2346 1886
rect 1362 1710 1372 1780
rect 1424 1710 1434 1780
rect 2287 1710 2293 1816
rect 2327 1710 2333 1816
rect 1375 1698 1421 1710
rect 2287 1698 2333 1710
rect 2429 1657 2604 1939
rect 2665 1886 2711 1898
rect 3577 1886 3623 1898
rect 2665 1780 2671 1886
rect 2705 1780 2711 1886
rect 3564 1816 3574 1886
rect 3626 1816 3636 1886
rect 2652 1710 2662 1780
rect 2714 1710 2724 1780
rect 3577 1710 3583 1816
rect 3617 1710 3623 1816
rect 2665 1698 2711 1710
rect 3577 1698 3623 1710
rect 3711 1657 3886 1939
rect 3955 1886 4001 1898
rect 4213 1886 4259 1898
rect 3955 1780 3961 1886
rect 3995 1780 4001 1886
rect 4200 1816 4210 1886
rect 4262 1816 4272 1886
rect 3942 1710 3952 1780
rect 4004 1710 4014 1780
rect 4213 1710 4219 1816
rect 4253 1710 4259 1816
rect 3955 1698 4001 1710
rect 4213 1698 4259 1710
rect 4304 1657 4418 1939
rect 4458 1902 4530 1910
rect 4458 1710 4468 1902
rect 4520 1710 4530 1902
rect 4471 1698 4517 1710
rect -495 1651 4461 1657
rect -495 1617 -225 1651
rect 63 1617 1065 1651
rect 1353 1617 2355 1651
rect 2643 1617 3645 1651
rect 3933 1617 4281 1651
rect 4449 1617 4461 1651
rect -495 1611 4461 1617
rect -633 1183 591 1189
rect -633 1149 -621 1183
rect -453 1149 -363 1183
rect -195 1149 -105 1183
rect 63 1149 153 1183
rect 321 1149 411 1183
rect 579 1149 591 1183
rect -633 1143 591 1149
rect 657 1183 1881 1189
rect 657 1149 669 1183
rect 837 1149 927 1183
rect 1095 1149 1185 1183
rect 1353 1149 1443 1183
rect 1611 1149 1701 1183
rect 1869 1149 1881 1183
rect 657 1143 1881 1149
rect 1947 1183 3171 1189
rect 1947 1149 1959 1183
rect 2127 1149 2217 1183
rect 2385 1149 2475 1183
rect 2643 1149 2733 1183
rect 2901 1149 2991 1183
rect 3159 1149 3171 1183
rect 1947 1143 3171 1149
rect 3237 1183 4461 1189
rect 3237 1149 3249 1183
rect 3417 1149 3507 1183
rect 3675 1149 3765 1183
rect 3933 1149 4023 1183
rect 4191 1149 4281 1183
rect 4449 1149 4461 1183
rect 3237 1143 4461 1149
rect -689 1099 -643 1111
rect -689 983 -683 1099
rect -649 983 -643 1099
rect -702 923 -692 983
rect -640 923 -630 983
rect -689 911 -643 923
rect -572 879 -505 1143
rect -431 1099 -385 1111
rect -431 983 -425 1099
rect -391 983 -385 1099
rect -444 923 -434 983
rect -382 923 -372 983
rect -431 911 -385 923
rect -314 879 -247 1143
rect -186 1099 -114 1143
rect -186 1039 -176 1099
rect -124 1039 -114 1099
rect -173 923 -167 1039
rect -133 923 -127 1039
rect -173 879 -127 923
rect -52 879 15 1143
rect 85 1099 131 1111
rect 85 983 91 1099
rect 125 983 131 1099
rect 72 923 82 983
rect 134 923 144 983
rect 85 911 131 923
rect 205 879 272 1143
rect 330 1099 402 1143
rect 330 1039 340 1099
rect 392 1039 402 1099
rect 343 923 349 1039
rect 383 923 389 1039
rect 343 879 389 923
rect 465 879 532 1143
rect 601 1099 647 1111
rect 601 983 607 1099
rect 641 983 647 1099
rect 588 923 598 983
rect 650 923 660 983
rect 601 911 647 923
rect 717 879 784 1143
rect 859 1099 905 1111
rect 859 983 865 1099
rect 899 983 905 1099
rect 846 923 856 983
rect 908 923 918 983
rect 859 911 905 923
rect 971 879 1038 1143
rect 1104 1099 1176 1143
rect 1104 1039 1114 1099
rect 1166 1039 1176 1099
rect 1117 923 1123 1039
rect 1157 923 1163 1039
rect 1117 879 1163 923
rect 1232 879 1299 1143
rect 1375 1099 1421 1111
rect 1375 983 1381 1099
rect 1415 983 1421 1099
rect 1362 923 1372 983
rect 1424 923 1434 983
rect 1375 911 1421 923
rect 1485 879 1552 1143
rect 1620 1099 1692 1143
rect 1620 1039 1630 1099
rect 1682 1039 1692 1099
rect 1633 923 1639 1039
rect 1673 923 1679 1039
rect 1633 879 1679 923
rect 1747 879 1814 1143
rect 1891 1099 1937 1111
rect 1891 983 1897 1099
rect 1931 983 1937 1099
rect 1878 923 1888 983
rect 1940 923 1950 983
rect 1891 911 1937 923
rect 2005 879 2072 1143
rect 2149 1099 2195 1111
rect 2149 983 2155 1099
rect 2189 983 2195 1099
rect 2136 923 2146 983
rect 2198 923 2208 983
rect 2149 911 2195 923
rect 2262 879 2329 1143
rect 2394 1099 2466 1143
rect 2394 1039 2404 1099
rect 2456 1039 2466 1099
rect 2407 923 2413 1039
rect 2447 923 2453 1039
rect 2407 879 2453 923
rect 2523 879 2590 1143
rect 2665 1099 2711 1111
rect 2665 983 2671 1099
rect 2705 983 2711 1099
rect 2652 923 2662 983
rect 2714 923 2724 983
rect 2665 911 2711 923
rect 2782 879 2849 1143
rect 2910 1099 2982 1143
rect 2910 1039 2920 1099
rect 2972 1039 2982 1099
rect 2923 923 2929 1039
rect 2963 923 2969 1039
rect 2923 879 2969 923
rect 3032 879 3099 1143
rect 3181 1099 3227 1111
rect 3181 983 3187 1099
rect 3221 983 3227 1099
rect 3168 923 3178 983
rect 3230 923 3240 983
rect 3181 911 3227 923
rect 3292 879 3359 1143
rect 3439 1099 3485 1111
rect 3439 983 3445 1099
rect 3479 983 3485 1099
rect 3426 923 3436 983
rect 3488 923 3498 983
rect 3439 911 3485 923
rect 3554 879 3621 1143
rect 3684 1099 3756 1143
rect 3684 1039 3694 1099
rect 3746 1039 3756 1099
rect 3697 923 3703 1039
rect 3737 923 3743 1039
rect 3697 879 3743 923
rect 3814 879 3881 1143
rect 3955 1099 4001 1111
rect 3955 983 3961 1099
rect 3995 983 4001 1099
rect 3942 923 3952 983
rect 4004 923 4014 983
rect 3955 911 4001 923
rect 4073 879 4140 1143
rect 4200 1099 4272 1143
rect 4200 1039 4210 1099
rect 4262 1039 4272 1099
rect 4213 923 4219 1039
rect 4253 923 4259 1039
rect 4213 879 4259 923
rect 4340 879 4407 1143
rect 4471 1099 4517 1111
rect 4458 1039 4468 1099
rect 4520 1039 4530 1099
rect 4471 983 4477 1039
rect 4511 983 4517 1039
rect 4458 923 4468 983
rect 4520 923 4530 983
rect 4471 911 4517 923
rect -633 873 591 879
rect -633 839 -621 873
rect -453 839 -363 873
rect -195 839 -105 873
rect 63 839 153 873
rect 321 839 411 873
rect 579 839 591 873
rect -633 833 591 839
rect 657 873 1881 879
rect 657 839 669 873
rect 837 839 927 873
rect 1095 839 1185 873
rect 1353 839 1443 873
rect 1611 839 1701 873
rect 1869 839 1881 873
rect 657 833 1881 839
rect 1947 873 3171 879
rect 1947 839 1959 873
rect 2127 839 2217 873
rect 2385 839 2475 873
rect 2643 839 2733 873
rect 2901 839 2991 873
rect 3159 839 3171 873
rect 1947 833 3171 839
rect 3237 873 4461 879
rect 3237 839 3249 873
rect 3417 839 3507 873
rect 3675 839 3765 873
rect 3933 839 4023 873
rect 4191 839 4281 873
rect 4449 839 4461 873
rect 3237 833 4461 839
rect -816 754 4615 760
rect -816 563 -804 754
rect 4603 563 4615 754
rect -816 557 4615 563
<< via1 >>
rect -374 2157 4658 2296
rect -296 1826 -287 1886
rect -287 1826 -253 1886
rect -253 1826 -244 1886
rect 994 1816 1003 1886
rect 1003 1816 1037 1886
rect 1037 1816 1046 1886
rect 82 1710 91 1770
rect 91 1710 125 1770
rect 125 1710 134 1770
rect 2284 1816 2293 1886
rect 2293 1816 2327 1886
rect 2327 1816 2336 1886
rect 1372 1710 1381 1780
rect 1381 1710 1415 1780
rect 1415 1710 1424 1780
rect 3574 1816 3583 1886
rect 3583 1816 3617 1886
rect 3617 1816 3626 1886
rect 2662 1710 2671 1780
rect 2671 1710 2705 1780
rect 2705 1710 2714 1780
rect 4210 1816 4219 1886
rect 4219 1816 4253 1886
rect 4253 1816 4262 1886
rect 3952 1710 3961 1780
rect 3961 1710 3995 1780
rect 3995 1710 4004 1780
rect 4468 1886 4520 1902
rect 4468 1710 4477 1886
rect 4477 1710 4511 1886
rect 4511 1710 4520 1886
rect -692 923 -683 983
rect -683 923 -649 983
rect -649 923 -640 983
rect -434 923 -425 983
rect -425 923 -391 983
rect -391 923 -382 983
rect -176 1039 -167 1099
rect -167 1039 -133 1099
rect -133 1039 -124 1099
rect 82 923 91 983
rect 91 923 125 983
rect 125 923 134 983
rect 340 1039 349 1099
rect 349 1039 383 1099
rect 383 1039 392 1099
rect 598 923 607 983
rect 607 923 641 983
rect 641 923 650 983
rect 856 923 865 983
rect 865 923 899 983
rect 899 923 908 983
rect 1114 1039 1123 1099
rect 1123 1039 1157 1099
rect 1157 1039 1166 1099
rect 1372 923 1381 983
rect 1381 923 1415 983
rect 1415 923 1424 983
rect 1630 1039 1639 1099
rect 1639 1039 1673 1099
rect 1673 1039 1682 1099
rect 1888 923 1897 983
rect 1897 923 1931 983
rect 1931 923 1940 983
rect 2146 923 2155 983
rect 2155 923 2189 983
rect 2189 923 2198 983
rect 2404 1039 2413 1099
rect 2413 1039 2447 1099
rect 2447 1039 2456 1099
rect 2662 923 2671 983
rect 2671 923 2705 983
rect 2705 923 2714 983
rect 2920 1039 2929 1099
rect 2929 1039 2963 1099
rect 2963 1039 2972 1099
rect 3178 923 3187 983
rect 3187 923 3221 983
rect 3221 923 3230 983
rect 3436 923 3445 983
rect 3445 923 3479 983
rect 3479 923 3488 983
rect 3694 1039 3703 1099
rect 3703 1039 3737 1099
rect 3737 1039 3746 1099
rect 3952 923 3961 983
rect 3961 923 3995 983
rect 3995 923 4004 983
rect 4210 1039 4219 1099
rect 4219 1039 4253 1099
rect 4253 1039 4262 1099
rect 4468 1039 4477 1099
rect 4477 1039 4511 1099
rect 4511 1039 4520 1099
rect 4468 923 4477 983
rect 4477 923 4511 983
rect 4511 923 4520 983
rect -804 563 4603 754
<< metal2 >>
rect -423 2296 4658 2306
rect -423 2157 -374 2296
rect -423 2147 4658 2157
rect -296 1886 -244 2147
rect -296 1816 -244 1826
rect 994 1886 1046 2147
rect 994 1806 1046 1816
rect 2284 1886 2336 2147
rect 2284 1806 2336 1816
rect 3574 1886 3626 2147
rect 3574 1806 3626 1816
rect 4210 1886 4262 2147
rect 4210 1806 4262 1816
rect 4468 1902 4520 1921
rect 1372 1780 1424 1790
rect 82 1770 134 1780
rect 82 1109 134 1710
rect 1372 1109 1424 1710
rect 2662 1780 2714 1790
rect 2662 1109 2714 1710
rect 3952 1780 4004 1790
rect 3952 1109 4004 1710
rect 4468 1474 4520 1710
rect 4468 1422 4746 1474
rect -176 1099 392 1109
rect -124 1039 340 1099
rect -176 1029 392 1039
rect 1114 1099 1682 1109
rect 1166 1039 1630 1099
rect 1114 1029 1682 1039
rect 2404 1099 2972 1109
rect 2456 1039 2920 1099
rect 2404 1029 2972 1039
rect 3694 1099 4262 1109
rect 3746 1039 4210 1099
rect 3694 1029 4262 1039
rect 4468 1099 4520 1422
rect 4468 993 4520 1039
rect -928 983 -640 993
rect -928 923 -692 983
rect -928 913 -640 923
rect -434 983 650 993
rect -382 923 82 983
rect 134 923 598 983
rect -434 913 650 923
rect 856 983 1940 993
rect 908 923 1372 983
rect 1424 923 1888 983
rect 856 913 1940 923
rect 2146 983 3230 993
rect 2198 923 2662 983
rect 2714 923 3178 983
rect 2146 913 3230 923
rect 3436 983 4520 993
rect 3488 923 3952 983
rect 4004 923 4468 983
rect 3436 913 4520 923
rect -897 754 4603 764
rect -897 563 -804 754
rect -897 553 4603 563
<< labels >>
rlabel metal2 -422 2228 -422 2228 3 vcc
port 1 e
rlabel metal2 4745 1450 4745 1450 3 vref
port 3 e
rlabel metal2 -896 637 -896 637 3 vss
port 2 e
rlabel metal2 -927 957 -927 957 3 vref0
port 4 e
rlabel metal1 -494 1637 -494 1637 3 vr
port 5 e
<< end >>
