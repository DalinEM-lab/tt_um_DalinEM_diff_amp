magic
tech sky130A
timestamp 1740708554
<< end >>
