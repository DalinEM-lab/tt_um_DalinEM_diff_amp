VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DalinEM_diff_amp
  CLASS BLOCK ;
  FOREIGN tt_um_DalinEM_diff_amp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.524000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 144.000000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 144.000000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 15.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 157.000 5.000 159.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.000 5.000 4.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 108.880 26.560 148.930 33.935 ;
      LAYER pwell ;
        RECT 108.900 8.990 114.000 15.950 ;
        RECT 115.200 6.335 142.835 24.110 ;
        RECT 115.620 6.165 115.735 6.335 ;
        RECT 116.205 6.165 142.370 6.175 ;
      LAYER li1 ;
        RECT 108.350 32.865 149.230 34.555 ;
        RECT 108.350 27.020 109.620 32.865 ;
        RECT 110.825 32.420 128.825 32.590 ;
        RECT 129.115 32.420 147.115 32.590 ;
        RECT 110.595 30.365 110.765 32.205 ;
        RECT 128.885 30.365 129.055 32.205 ;
        RECT 147.175 30.365 147.345 32.205 ;
        RECT 110.825 29.980 128.825 30.150 ;
        RECT 129.115 29.980 147.115 30.150 ;
        RECT 110.595 27.925 110.765 29.765 ;
        RECT 128.885 27.925 129.055 29.765 ;
        RECT 147.175 27.925 147.345 29.765 ;
        RECT 110.825 27.540 128.825 27.710 ;
        RECT 129.115 27.540 147.115 27.710 ;
        RECT 148.180 27.020 149.225 32.865 ;
        RECT 108.350 26.355 149.225 27.020 ;
        RECT 108.355 23.480 144.100 24.180 ;
        RECT 108.355 15.775 115.735 23.480 ;
        RECT 116.875 23.015 128.875 23.185 ;
        RECT 129.165 23.015 141.165 23.185 ;
        RECT 116.645 16.805 116.815 22.845 ;
        RECT 128.935 16.805 129.105 22.845 ;
        RECT 141.225 16.805 141.395 22.845 ;
        RECT 116.875 16.465 128.875 16.635 ;
        RECT 129.165 16.465 141.165 16.635 ;
        RECT 108.350 15.590 115.735 15.775 ;
        RECT 108.350 9.360 109.405 15.590 ;
        RECT 109.930 15.030 112.970 15.200 ;
        RECT 109.590 9.970 109.760 14.970 ;
        RECT 113.140 9.970 113.310 14.970 ;
        RECT 109.930 9.360 112.970 9.910 ;
        RECT 113.610 9.360 115.735 15.590 ;
        RECT 116.870 13.640 128.870 13.810 ;
        RECT 129.160 13.640 141.160 13.810 ;
        RECT 108.350 8.210 115.735 9.360 ;
        RECT 108.340 6.810 115.735 8.210 ;
        RECT 116.640 7.430 116.810 13.470 ;
        RECT 128.930 7.430 129.100 13.470 ;
        RECT 141.220 7.430 141.390 13.470 ;
        RECT 116.870 7.090 128.870 7.260 ;
        RECT 129.160 7.090 141.160 7.260 ;
        RECT 142.350 6.810 144.100 23.480 ;
        RECT 108.340 5.260 144.100 6.810 ;
      LAYER met1 ;
        RECT 109.210 33.900 148.320 34.405 ;
        RECT 109.860 32.390 147.095 32.620 ;
        RECT 109.860 30.380 110.860 32.390 ;
        RECT 109.860 25.225 110.290 30.380 ;
        RECT 111.745 30.180 127.940 32.390 ;
        RECT 128.855 32.125 129.085 32.185 ;
        RECT 128.785 30.445 129.155 32.125 ;
        RECT 128.855 30.385 129.085 30.445 ;
        RECT 130.055 30.180 146.250 32.390 ;
        RECT 147.075 30.390 148.085 32.190 ;
        RECT 147.145 30.385 147.375 30.390 ;
        RECT 110.845 29.950 128.805 30.180 ;
        RECT 129.135 29.950 147.095 30.180 ;
        RECT 110.430 27.940 110.860 29.745 ;
        RECT 111.745 27.740 127.940 29.950 ;
        RECT 128.855 29.685 129.085 29.745 ;
        RECT 128.785 28.005 129.155 29.685 ;
        RECT 128.855 27.945 129.085 28.005 ;
        RECT 130.055 27.740 146.250 29.950 ;
        RECT 147.085 27.740 147.515 29.745 ;
        RECT 110.845 27.510 147.515 27.740 ;
        RECT 147.655 26.150 148.085 30.390 ;
        RECT 110.430 25.650 152.710 26.150 ;
        RECT 109.860 24.725 147.565 25.225 ;
        RECT 151.810 24.470 152.710 25.650 ;
        RECT 116.895 22.985 128.855 23.215 ;
        RECT 129.185 22.985 141.145 23.215 ;
        RECT 116.615 22.765 116.845 22.825 ;
        RECT 116.375 17.095 116.905 22.765 ;
        RECT 116.615 16.825 116.845 17.095 ;
        RECT 120.135 16.695 125.560 22.985 ;
        RECT 128.905 18.640 129.135 22.825 ;
        RECT 128.845 17.045 129.205 18.640 ;
        RECT 128.905 16.825 129.135 17.045 ;
        RECT 132.655 16.695 138.090 22.985 ;
        RECT 141.195 22.765 141.425 22.825 ;
        RECT 141.135 17.160 141.665 22.765 ;
        RECT 141.195 16.825 141.425 17.160 ;
        RECT 116.925 16.665 128.845 16.695 ;
        RECT 129.195 16.665 141.135 16.695 ;
        RECT 116.895 16.435 128.855 16.665 ;
        RECT 129.185 16.435 141.145 16.665 ;
        RECT 116.925 16.410 128.845 16.435 ;
        RECT 129.195 16.410 141.135 16.435 ;
        RECT 116.975 15.730 130.290 16.125 ;
        RECT 109.960 15.230 112.940 15.285 ;
        RECT 109.950 15.000 112.950 15.230 ;
        RECT 109.560 13.955 109.790 14.950 ;
        RECT 113.110 14.045 113.405 14.950 ;
        RECT 127.740 14.195 141.085 14.640 ;
        RECT 113.050 13.955 113.410 14.045 ;
        RECT 109.560 10.970 113.410 13.955 ;
        RECT 116.900 13.840 128.840 13.870 ;
        RECT 129.190 13.840 141.130 13.865 ;
        RECT 116.890 13.610 128.850 13.840 ;
        RECT 129.180 13.610 141.140 13.840 ;
        RECT 116.900 13.585 128.840 13.610 ;
        RECT 116.610 13.390 116.840 13.450 ;
        RECT 109.560 9.990 109.790 10.970 ;
        RECT 113.050 10.050 113.410 10.970 ;
        RECT 113.110 9.990 113.405 10.050 ;
        RECT 109.950 9.710 112.950 9.940 ;
        RECT 115.845 7.685 116.900 13.390 ;
        RECT 116.610 7.450 116.840 7.685 ;
        RECT 120.110 7.295 125.545 13.585 ;
        RECT 129.190 13.580 141.130 13.610 ;
        RECT 128.900 13.235 129.130 13.450 ;
        RECT 128.840 11.640 129.200 13.235 ;
        RECT 128.900 7.450 129.130 11.640 ;
        RECT 108.820 6.690 111.705 7.220 ;
        RECT 116.890 7.035 128.850 7.295 ;
        RECT 129.190 7.290 131.690 7.300 ;
        RECT 132.610 7.290 138.045 13.580 ;
        RECT 141.190 13.390 141.420 13.450 ;
        RECT 141.125 8.030 141.985 13.390 ;
        RECT 141.190 7.450 141.420 8.030 ;
        RECT 129.180 7.060 141.140 7.290 ;
        RECT 129.190 7.040 131.690 7.060 ;
        RECT 108.830 5.540 143.620 6.045 ;
      LAYER met2 ;
        RECT 108.350 33.885 154.395 35.880 ;
        RECT 108.350 33.880 151.230 33.885 ;
        RECT 110.380 26.165 110.810 29.745 ;
        RECT 128.835 27.955 129.105 33.880 ;
        RECT 110.380 25.645 111.975 26.165 ;
        RECT 114.470 25.650 116.275 26.150 ;
        RECT 139.790 25.650 141.615 26.150 ;
        RECT 110.010 14.960 112.890 15.385 ;
        RECT 113.100 14.090 113.360 14.095 ;
        RECT 113.085 10.000 113.375 14.090 ;
        RECT 115.845 13.440 116.275 25.650 ;
        RECT 116.425 24.725 118.355 25.225 ;
        RECT 116.425 19.875 116.855 24.725 ;
        RECT 141.185 19.875 141.615 25.650 ;
        RECT 147.135 25.225 147.565 29.745 ;
        RECT 141.765 24.725 143.635 25.225 ;
        RECT 145.460 24.725 147.565 25.225 ;
        RECT 128.875 16.945 129.155 18.755 ;
        RECT 116.975 15.770 118.025 16.745 ;
        RECT 127.740 13.535 128.790 14.580 ;
        RECT 129.240 13.530 130.290 16.185 ;
        RECT 140.035 14.205 141.085 16.745 ;
        RECT 141.765 13.440 142.195 24.725 ;
        RECT 151.860 24.420 152.660 26.150 ;
        RECT 115.845 10.570 116.850 13.440 ;
        RECT 128.870 11.540 129.160 13.335 ;
        RECT 115.845 7.685 116.860 10.570 ;
        RECT 141.175 7.980 142.195 13.440 ;
        RECT 108.340 7.515 112.250 7.520 ;
        RECT 66.720 6.065 112.250 7.515 ;
        RECT 116.950 6.970 119.350 7.360 ;
        RECT 129.240 6.980 131.640 7.370 ;
        RECT 66.720 5.520 143.560 6.065 ;
        RECT 66.720 5.515 89.070 5.520 ;
      LAYER met3 ;
        RECT 150.435 33.885 154.430 35.875 ;
        RECT 151.810 24.445 152.710 26.125 ;
        RECT 128.820 15.360 129.210 18.730 ;
        RECT 109.960 14.985 129.210 15.360 ;
        RECT 66.670 5.520 70.465 7.510 ;
        RECT 113.035 5.140 113.935 14.065 ;
        RECT 128.820 11.565 129.210 14.985 ;
        RECT 93.850 4.240 113.935 5.140 ;
        RECT 116.900 6.995 119.400 7.335 ;
        RECT 129.190 7.005 131.690 7.345 ;
        RECT 116.900 3.910 117.800 6.995 ;
        RECT 115.160 3.020 117.800 3.910 ;
        RECT 116.900 3.015 117.800 3.020 ;
        RECT 129.190 3.910 130.090 7.005 ;
        RECT 129.190 3.020 131.870 3.910 ;
        RECT 129.190 3.015 130.090 3.020 ;
      LAYER met4 ;
        RECT 30.670 220.760 30.970 224.760 ;
        RECT 33.430 220.760 33.730 224.760 ;
        RECT 36.190 220.760 36.490 224.760 ;
        RECT 38.950 220.760 39.250 224.760 ;
        RECT 41.710 220.760 42.010 224.760 ;
        RECT 44.470 220.760 44.770 224.760 ;
        RECT 47.230 220.760 47.530 224.760 ;
        RECT 49.990 220.760 50.290 224.760 ;
        RECT 52.750 220.760 53.050 224.760 ;
        RECT 55.510 220.760 55.810 224.760 ;
        RECT 58.270 220.760 58.570 224.760 ;
        RECT 61.030 220.760 61.330 224.760 ;
        RECT 63.790 220.760 64.090 224.760 ;
        RECT 66.550 220.760 66.850 224.760 ;
        RECT 69.310 220.760 69.610 224.760 ;
        RECT 72.070 220.760 72.370 224.760 ;
        RECT 74.830 220.760 75.130 224.760 ;
        RECT 77.590 220.760 77.890 224.760 ;
        RECT 80.350 220.760 80.650 224.760 ;
        RECT 83.110 220.760 83.410 224.760 ;
        RECT 85.870 220.760 86.170 224.760 ;
        RECT 88.630 220.760 88.930 224.760 ;
        RECT 91.390 220.760 91.690 224.760 ;
        RECT 94.150 220.760 94.450 224.760 ;
        RECT 4.000 218.760 94.450 220.760 ;
        RECT 150.025 33.880 157.000 35.880 ;
        RECT 4.000 5.515 70.420 7.515 ;
        RECT 93.850 4.240 96.385 5.140 ;
        RECT 93.850 1.000 94.750 4.240 ;
        RECT 113.170 3.015 117.800 3.915 ;
        RECT 129.190 3.015 133.390 3.915 ;
        RECT 113.170 1.000 114.070 3.015 ;
        RECT 132.490 1.000 133.390 3.015 ;
        RECT 151.810 1.000 152.710 26.150 ;
  END
END tt_um_DalinEM_diff_amp
END LIBRARY

