magic
tech sky130A
magscale 1 2
timestamp 1741058913
<< metal3 >>
rect -1886 1712 1886 1740
rect -1886 -1712 1802 1712
rect 1866 -1712 1886 1712
rect -1886 -1740 1886 -1712
<< via3 >>
rect 1802 -1712 1866 1712
<< mimcap >>
rect -1846 1660 1554 1700
rect -1846 -1660 -1806 1660
rect 1514 -1660 1554 1660
rect -1846 -1700 1554 -1660
<< mimcapcontact >>
rect -1806 -1660 1514 1660
<< metal4 >>
rect 1786 1712 1882 1728
rect -1807 1660 1515 1661
rect -1807 -1660 -1806 1660
rect 1514 -1660 1515 1660
rect -1807 -1661 1515 -1660
rect 1786 -1712 1802 1712
rect 1866 -1712 1882 1712
rect 1786 -1728 1882 -1712
<< properties >>
string FIXED_BBOX -1886 -1740 1594 1740
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17.0 l 17.0 val 590.92 carea 2.00 cperi 0.19 class capacitor nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100 mf 1
<< end >>
