VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DalinEM_diff_amp
  CLASS BLOCK ;
  FOREIGN tt_um_DalinEM_diff_amp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.524000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 144.000000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 144.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 15.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.595499 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 157.000 5.000 159.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.000 5.000 4.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 89.560 26.555 129.610 33.930 ;
      LAYER pwell ;
        RECT 89.580 8.985 94.680 15.945 ;
        RECT 95.880 6.330 123.515 24.105 ;
        RECT 96.300 6.160 96.415 6.330 ;
        RECT 96.885 6.160 123.050 6.170 ;
      LAYER li1 ;
        RECT 89.030 32.860 129.910 34.550 ;
        RECT 89.030 27.015 90.300 32.860 ;
        RECT 91.505 32.415 109.505 32.585 ;
        RECT 109.795 32.415 127.795 32.585 ;
        RECT 91.275 30.360 91.445 32.200 ;
        RECT 109.565 30.360 109.735 32.200 ;
        RECT 127.855 30.360 128.025 32.200 ;
        RECT 91.505 29.975 109.505 30.145 ;
        RECT 109.795 29.975 127.795 30.145 ;
        RECT 91.275 27.920 91.445 29.760 ;
        RECT 109.565 27.920 109.735 29.760 ;
        RECT 127.855 27.920 128.025 29.760 ;
        RECT 91.505 27.535 109.505 27.705 ;
        RECT 109.795 27.535 127.795 27.705 ;
        RECT 128.860 27.015 129.905 32.860 ;
        RECT 89.030 26.350 129.905 27.015 ;
        RECT 89.035 23.475 124.780 24.175 ;
        RECT 89.035 15.770 96.415 23.475 ;
        RECT 97.555 23.010 109.555 23.180 ;
        RECT 109.845 23.010 121.845 23.180 ;
        RECT 97.325 16.800 97.495 22.840 ;
        RECT 109.615 16.800 109.785 22.840 ;
        RECT 121.905 16.800 122.075 22.840 ;
        RECT 97.555 16.460 109.555 16.630 ;
        RECT 109.845 16.460 121.845 16.630 ;
        RECT 89.030 15.585 96.415 15.770 ;
        RECT 89.030 9.355 90.085 15.585 ;
        RECT 90.610 15.025 93.650 15.195 ;
        RECT 90.270 9.965 90.440 14.965 ;
        RECT 93.820 9.965 93.990 14.965 ;
        RECT 90.610 9.355 93.650 9.905 ;
        RECT 94.290 9.355 96.415 15.585 ;
        RECT 97.550 13.635 109.550 13.805 ;
        RECT 109.840 13.635 121.840 13.805 ;
        RECT 89.030 8.205 96.415 9.355 ;
        RECT 89.020 6.805 96.415 8.205 ;
        RECT 97.320 7.425 97.490 13.465 ;
        RECT 109.610 7.425 109.780 13.465 ;
        RECT 121.900 7.425 122.070 13.465 ;
        RECT 97.550 7.085 109.550 7.255 ;
        RECT 109.840 7.085 121.840 7.255 ;
        RECT 123.030 6.805 124.780 23.475 ;
        RECT 89.020 5.255 124.780 6.805 ;
      LAYER met1 ;
        RECT 89.890 33.895 129.000 34.400 ;
        RECT 90.540 32.385 127.775 32.615 ;
        RECT 90.540 30.375 91.540 32.385 ;
        RECT 90.540 25.220 90.970 30.375 ;
        RECT 92.425 30.175 108.620 32.385 ;
        RECT 109.535 32.120 109.765 32.180 ;
        RECT 109.465 30.440 109.835 32.120 ;
        RECT 109.535 30.380 109.765 30.440 ;
        RECT 110.735 30.175 126.930 32.385 ;
        RECT 127.755 30.385 128.765 32.185 ;
        RECT 127.825 30.380 128.055 30.385 ;
        RECT 91.525 29.945 109.485 30.175 ;
        RECT 109.815 29.945 127.775 30.175 ;
        RECT 91.110 27.935 91.540 29.740 ;
        RECT 92.425 27.735 108.620 29.945 ;
        RECT 109.535 29.680 109.765 29.740 ;
        RECT 109.465 28.000 109.835 29.680 ;
        RECT 109.535 27.940 109.765 28.000 ;
        RECT 110.735 27.735 126.930 29.945 ;
        RECT 127.765 27.735 128.195 29.740 ;
        RECT 91.525 27.505 128.195 27.735 ;
        RECT 128.335 26.145 128.765 30.385 ;
        RECT 91.110 25.645 133.390 26.145 ;
        RECT 90.540 24.720 128.245 25.220 ;
        RECT 132.490 24.465 133.390 25.645 ;
        RECT 97.575 22.980 109.535 23.210 ;
        RECT 109.865 22.980 121.825 23.210 ;
        RECT 97.295 22.760 97.525 22.820 ;
        RECT 97.055 17.090 97.585 22.760 ;
        RECT 97.295 16.820 97.525 17.090 ;
        RECT 100.815 16.690 106.240 22.980 ;
        RECT 109.585 18.635 109.815 22.820 ;
        RECT 109.525 17.040 109.885 18.635 ;
        RECT 109.585 16.820 109.815 17.040 ;
        RECT 113.335 16.690 118.770 22.980 ;
        RECT 121.875 22.760 122.105 22.820 ;
        RECT 121.815 17.155 122.345 22.760 ;
        RECT 121.875 16.820 122.105 17.155 ;
        RECT 97.605 16.660 109.525 16.690 ;
        RECT 109.875 16.660 121.815 16.690 ;
        RECT 97.575 16.430 109.535 16.660 ;
        RECT 109.865 16.430 121.825 16.660 ;
        RECT 97.605 16.405 109.525 16.430 ;
        RECT 109.875 16.405 121.815 16.430 ;
        RECT 97.655 15.725 110.970 16.120 ;
        RECT 90.640 15.225 93.620 15.280 ;
        RECT 90.630 14.995 93.630 15.225 ;
        RECT 90.240 13.950 90.470 14.945 ;
        RECT 93.790 14.040 94.085 14.945 ;
        RECT 108.420 14.190 121.765 14.635 ;
        RECT 93.730 13.950 94.090 14.040 ;
        RECT 90.240 10.965 94.090 13.950 ;
        RECT 97.580 13.835 109.520 13.865 ;
        RECT 109.870 13.835 121.810 13.860 ;
        RECT 97.570 13.605 109.530 13.835 ;
        RECT 109.860 13.605 121.820 13.835 ;
        RECT 97.580 13.580 109.520 13.605 ;
        RECT 97.290 13.385 97.520 13.445 ;
        RECT 90.240 9.985 90.470 10.965 ;
        RECT 93.730 10.045 94.090 10.965 ;
        RECT 93.790 9.985 94.085 10.045 ;
        RECT 90.630 9.705 93.630 9.935 ;
        RECT 96.525 7.680 97.580 13.385 ;
        RECT 97.290 7.445 97.520 7.680 ;
        RECT 100.790 7.290 106.225 13.580 ;
        RECT 109.870 13.575 121.810 13.605 ;
        RECT 109.580 13.230 109.810 13.445 ;
        RECT 109.520 11.635 109.880 13.230 ;
        RECT 109.580 7.445 109.810 11.635 ;
        RECT 89.500 6.685 92.385 7.215 ;
        RECT 97.570 7.030 109.530 7.290 ;
        RECT 109.870 7.285 112.370 7.295 ;
        RECT 113.290 7.285 118.725 13.575 ;
        RECT 121.870 13.385 122.100 13.445 ;
        RECT 121.805 8.025 122.665 13.385 ;
        RECT 121.870 7.445 122.100 8.025 ;
        RECT 109.860 7.055 121.820 7.285 ;
        RECT 109.870 7.035 112.370 7.055 ;
        RECT 89.510 5.535 124.300 6.040 ;
      LAYER met2 ;
        RECT 89.030 33.880 134.275 35.875 ;
        RECT 89.030 33.875 131.110 33.880 ;
        RECT 91.060 26.160 91.490 29.740 ;
        RECT 109.515 27.950 109.785 33.875 ;
        RECT 91.060 25.640 92.655 26.160 ;
        RECT 95.150 25.645 96.955 26.145 ;
        RECT 120.470 25.645 122.295 26.145 ;
        RECT 90.690 14.955 93.570 15.380 ;
        RECT 93.780 14.085 94.040 14.090 ;
        RECT 93.765 9.995 94.055 14.085 ;
        RECT 96.525 13.435 96.955 25.645 ;
        RECT 97.105 24.720 99.035 25.220 ;
        RECT 97.105 19.870 97.535 24.720 ;
        RECT 121.865 19.870 122.295 25.645 ;
        RECT 127.815 25.220 128.245 29.740 ;
        RECT 122.445 24.720 124.315 25.220 ;
        RECT 126.140 24.720 128.245 25.220 ;
        RECT 109.555 16.940 109.835 18.750 ;
        RECT 97.655 15.765 98.705 16.740 ;
        RECT 108.420 13.530 109.470 14.575 ;
        RECT 109.920 13.525 110.970 16.180 ;
        RECT 120.715 14.200 121.765 16.740 ;
        RECT 122.445 13.435 122.875 24.720 ;
        RECT 132.540 24.415 133.340 26.145 ;
        RECT 96.525 10.565 97.530 13.435 ;
        RECT 109.550 11.535 109.840 13.330 ;
        RECT 96.525 7.680 97.540 10.565 ;
        RECT 121.855 7.975 122.875 13.435 ;
        RECT 66.720 6.060 92.930 7.515 ;
        RECT 97.630 6.965 100.030 7.355 ;
        RECT 109.920 6.975 112.320 7.365 ;
        RECT 66.720 5.515 124.240 6.060 ;
      LAYER met3 ;
        RECT 130.315 33.880 134.325 35.870 ;
        RECT 132.490 24.440 133.390 26.120 ;
        RECT 109.500 15.355 109.890 18.725 ;
        RECT 90.640 14.980 109.890 15.355 ;
        RECT 66.670 5.520 70.465 7.510 ;
        RECT 93.715 5.140 94.615 14.060 ;
        RECT 109.500 11.560 109.890 14.980 ;
        RECT 74.530 4.240 94.615 5.140 ;
        RECT 97.580 6.990 100.080 7.330 ;
        RECT 109.870 7.000 112.370 7.340 ;
        RECT 97.580 3.910 98.480 6.990 ;
        RECT 95.840 3.020 98.480 3.910 ;
        RECT 97.580 3.015 98.480 3.020 ;
        RECT 109.870 3.910 110.770 7.000 ;
        RECT 109.870 3.020 112.550 3.910 ;
        RECT 109.870 3.015 110.770 3.020 ;
      LAYER met4 ;
        RECT 30.670 220.760 30.970 224.760 ;
        RECT 33.430 220.760 33.730 224.760 ;
        RECT 36.190 220.760 36.490 224.760 ;
        RECT 38.950 220.760 39.250 224.760 ;
        RECT 41.710 220.760 42.010 224.760 ;
        RECT 44.470 220.760 44.770 224.760 ;
        RECT 47.230 220.760 47.530 224.760 ;
        RECT 49.990 220.760 50.290 224.760 ;
        RECT 52.750 220.760 53.050 224.760 ;
        RECT 55.510 220.760 55.810 224.760 ;
        RECT 58.270 220.760 58.570 224.760 ;
        RECT 61.030 220.760 61.330 224.760 ;
        RECT 63.790 220.760 64.090 224.760 ;
        RECT 66.550 220.760 66.850 224.760 ;
        RECT 69.310 220.760 69.610 224.760 ;
        RECT 72.070 220.760 72.370 224.760 ;
        RECT 74.830 220.760 75.130 224.760 ;
        RECT 77.590 220.760 77.890 224.760 ;
        RECT 80.350 220.760 80.650 224.760 ;
        RECT 83.110 220.760 83.410 224.760 ;
        RECT 85.870 220.760 86.170 224.760 ;
        RECT 88.630 220.760 88.930 224.760 ;
        RECT 91.390 220.760 91.690 224.760 ;
        RECT 94.150 220.760 94.450 224.760 ;
        RECT 4.000 218.760 94.450 220.760 ;
        RECT 129.905 33.875 157.000 35.875 ;
        RECT 4.000 5.515 70.420 7.515 ;
        RECT 74.530 4.240 77.065 5.140 ;
        RECT 74.530 1.000 75.430 4.240 ;
        RECT 93.850 3.015 98.480 3.915 ;
        RECT 109.870 3.015 114.070 3.915 ;
        RECT 93.850 1.000 94.750 3.015 ;
        RECT 113.170 1.000 114.070 3.015 ;
        RECT 132.490 1.000 133.390 26.145 ;
  END
END tt_um_DalinEM_diff_amp
END LIBRARY

