VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DalinEM_diff_amp
  CLASS BLOCK ;
  FOREIGN tt_um_DalinEM_diff_amp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.044000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.524000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 288.000000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 288.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 15.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 53.457798 ;
    ANTENNADIFFAREA 185.774292 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 157.005 5.000 159.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.000 5.000 4.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 16.615 146.635 56.665 154.010 ;
      LAYER pwell ;
        RECT 16.635 129.065 21.735 136.025 ;
        RECT 22.935 126.410 50.570 144.185 ;
        RECT 23.355 126.240 23.470 126.410 ;
        RECT 23.940 126.240 50.105 126.250 ;
      LAYER nwell ;
        RECT 58.905 126.245 71.970 165.040 ;
        RECT 84.085 126.890 94.115 136.080 ;
        RECT 103.715 127.340 128.185 139.510 ;
      LAYER pwell ;
        RECT 110.595 115.240 121.275 126.665 ;
      LAYER nwell ;
        RECT 126.215 121.190 130.305 125.980 ;
      LAYER pwell ;
        RECT 60.250 86.080 75.820 109.330 ;
        RECT 60.250 85.920 66.470 86.080 ;
        RECT 66.490 86.075 75.820 86.080 ;
        RECT 66.490 85.920 66.720 86.075 ;
        RECT 60.250 85.910 66.720 85.920 ;
        RECT 66.735 85.910 75.820 86.075 ;
        RECT 60.250 75.120 75.820 85.910 ;
        RECT 78.800 84.680 83.035 113.050 ;
      LAYER nwell ;
        RECT 83.340 106.115 86.515 112.980 ;
      LAYER pwell ;
        RECT 112.220 109.250 119.820 114.500 ;
        RECT 123.615 113.900 130.635 115.910 ;
      LAYER nwell ;
        RECT 83.260 99.635 86.450 103.595 ;
        RECT 83.260 93.185 86.450 97.145 ;
        RECT 83.260 86.735 86.450 90.695 ;
      LAYER pwell ;
        RECT 76.050 81.325 82.750 82.090 ;
        RECT 76.050 76.155 76.815 81.325 ;
        RECT 81.985 76.155 82.750 81.325 ;
      LAYER nwell ;
        RECT 83.295 81.110 86.455 85.265 ;
      LAYER pwell ;
        RECT 76.050 75.390 82.750 76.155 ;
      LAYER nwell ;
        RECT 83.290 75.210 86.455 81.110 ;
        RECT 83.290 75.190 86.450 75.210 ;
      LAYER pwell ;
        RECT 13.425 41.735 28.995 52.525 ;
      LAYER nwell ;
        RECT 36.465 52.435 39.625 52.455 ;
      LAYER pwell ;
        RECT 29.225 51.490 35.925 52.255 ;
        RECT 29.225 46.320 29.990 51.490 ;
        RECT 35.160 46.320 35.925 51.490 ;
      LAYER nwell ;
        RECT 36.465 46.535 39.630 52.435 ;
        RECT 89.160 47.705 129.210 55.080 ;
      LAYER pwell ;
        RECT 29.225 45.555 35.925 46.320 ;
        RECT 13.425 41.725 19.895 41.735 ;
        RECT 13.425 41.565 19.645 41.725 ;
        RECT 19.665 41.570 19.895 41.725 ;
        RECT 19.910 41.570 28.995 41.735 ;
        RECT 19.665 41.565 28.995 41.570 ;
        RECT 13.425 18.315 28.995 41.565 ;
        RECT 31.975 14.100 36.210 42.470 ;
      LAYER nwell ;
        RECT 36.470 42.380 39.630 46.535 ;
        RECT 36.435 36.455 39.625 40.415 ;
        RECT 36.435 30.005 39.625 33.965 ;
      LAYER pwell ;
        RECT 89.180 30.135 94.280 37.095 ;
      LAYER nwell ;
        RECT 36.435 23.555 39.625 27.515 ;
      LAYER pwell ;
        RECT 95.480 27.480 123.115 45.255 ;
        RECT 95.900 27.310 96.015 27.480 ;
        RECT 96.485 27.310 122.650 27.320 ;
      LAYER nwell ;
        RECT 36.515 14.170 39.690 21.035 ;
      LAYER li1 ;
        RECT 58.830 163.955 72.155 165.125 ;
        RECT 16.085 152.940 56.965 154.630 ;
        RECT 16.085 147.095 17.355 152.940 ;
        RECT 18.560 152.495 36.560 152.665 ;
        RECT 36.850 152.495 54.850 152.665 ;
        RECT 18.330 150.440 18.500 152.280 ;
        RECT 36.620 150.440 36.790 152.280 ;
        RECT 54.910 150.440 55.080 152.280 ;
        RECT 18.560 150.055 36.560 150.225 ;
        RECT 36.850 150.055 54.850 150.225 ;
        RECT 18.330 148.000 18.500 149.840 ;
        RECT 36.620 148.000 36.790 149.840 ;
        RECT 54.910 148.000 55.080 149.840 ;
        RECT 18.560 147.615 36.560 147.785 ;
        RECT 36.850 147.615 54.850 147.785 ;
        RECT 55.915 147.095 56.960 152.940 ;
        RECT 16.085 146.430 56.960 147.095 ;
        RECT 16.090 143.555 51.835 144.255 ;
        RECT 16.090 135.850 23.470 143.555 ;
        RECT 24.610 143.090 36.610 143.260 ;
        RECT 36.900 143.090 48.900 143.260 ;
        RECT 24.380 136.880 24.550 142.920 ;
        RECT 36.670 136.880 36.840 142.920 ;
        RECT 48.960 136.880 49.130 142.920 ;
        RECT 24.610 136.540 36.610 136.710 ;
        RECT 36.900 136.540 48.900 136.710 ;
        RECT 16.085 135.665 23.470 135.850 ;
        RECT 16.085 129.435 17.140 135.665 ;
        RECT 17.665 135.105 20.705 135.275 ;
        RECT 17.325 130.045 17.495 135.045 ;
        RECT 20.875 130.045 21.045 135.045 ;
        RECT 17.665 129.435 20.705 129.985 ;
        RECT 21.345 129.435 23.470 135.665 ;
        RECT 24.605 133.715 36.605 133.885 ;
        RECT 36.895 133.715 48.895 133.885 ;
        RECT 16.085 128.285 23.470 129.435 ;
        RECT 16.075 126.885 23.470 128.285 ;
        RECT 24.375 127.505 24.545 133.545 ;
        RECT 36.665 127.505 36.835 133.545 ;
        RECT 48.955 127.505 49.125 133.545 ;
        RECT 24.605 127.165 36.605 127.335 ;
        RECT 36.895 127.165 48.895 127.335 ;
        RECT 50.085 126.885 51.835 143.555 ;
        RECT 16.075 125.335 51.835 126.885 ;
        RECT 58.830 126.940 60.000 163.955 ;
        RECT 60.920 162.875 62.820 163.045 ;
        RECT 63.110 162.875 65.010 163.045 ;
        RECT 65.300 162.875 67.200 163.045 ;
        RECT 67.490 162.875 69.390 163.045 ;
        RECT 60.690 147.620 60.860 162.660 ;
        RECT 62.880 147.620 63.050 162.660 ;
        RECT 65.070 147.620 65.240 162.660 ;
        RECT 67.260 147.620 67.430 162.660 ;
        RECT 69.450 147.620 69.620 162.660 ;
        RECT 60.920 147.235 62.820 147.405 ;
        RECT 63.110 147.235 65.010 147.405 ;
        RECT 65.300 147.235 67.200 147.405 ;
        RECT 67.490 147.235 69.390 147.405 ;
        RECT 60.920 142.990 62.820 143.160 ;
        RECT 63.110 142.990 65.010 143.160 ;
        RECT 65.300 142.990 67.200 143.160 ;
        RECT 67.490 142.990 69.390 143.160 ;
        RECT 60.690 127.735 60.860 142.775 ;
        RECT 62.880 127.735 63.050 142.775 ;
        RECT 65.070 127.735 65.240 142.775 ;
        RECT 67.260 127.735 67.430 142.775 ;
        RECT 69.450 127.735 69.620 142.775 ;
        RECT 70.575 137.930 72.155 163.955 ;
        RECT 102.750 139.130 128.400 142.650 ;
        RECT 102.750 138.400 128.415 139.130 ;
        RECT 70.575 135.600 95.855 137.930 ;
        RECT 60.920 127.350 62.820 127.520 ;
        RECT 63.110 127.350 65.010 127.520 ;
        RECT 65.300 127.350 67.200 127.520 ;
        RECT 67.490 127.350 69.390 127.520 ;
        RECT 70.575 126.940 72.155 135.600 ;
        RECT 58.830 126.250 72.155 126.940 ;
        RECT 82.775 127.385 84.485 135.600 ;
        RECT 85.065 135.220 86.865 135.390 ;
        RECT 87.155 135.220 88.955 135.390 ;
        RECT 89.245 135.220 91.045 135.390 ;
        RECT 91.335 135.220 93.135 135.390 ;
        RECT 84.835 127.965 85.005 135.005 ;
        RECT 86.925 127.965 87.095 135.005 ;
        RECT 89.015 127.965 89.185 135.005 ;
        RECT 91.105 127.965 91.275 135.005 ;
        RECT 93.195 127.965 93.365 135.005 ;
        RECT 85.065 127.580 86.865 127.750 ;
        RECT 87.155 127.580 88.955 127.750 ;
        RECT 89.245 127.580 91.045 127.750 ;
        RECT 91.335 127.580 93.135 127.750 ;
        RECT 93.685 127.385 95.855 135.600 ;
        RECT 82.775 127.285 95.855 127.385 ;
        RECT 103.705 128.120 104.605 138.400 ;
        RECT 105.530 137.945 110.530 138.115 ;
        RECT 110.820 137.945 115.820 138.115 ;
        RECT 116.110 137.945 121.110 138.115 ;
        RECT 121.400 137.945 126.400 138.115 ;
        RECT 105.300 135.190 105.470 137.730 ;
        RECT 110.590 135.190 110.760 137.730 ;
        RECT 115.880 135.190 116.050 137.730 ;
        RECT 121.170 135.190 121.340 137.730 ;
        RECT 126.460 135.190 126.630 137.730 ;
        RECT 105.530 134.805 110.530 134.975 ;
        RECT 110.820 134.805 115.820 134.975 ;
        RECT 116.110 134.805 121.110 134.975 ;
        RECT 121.400 134.805 126.400 134.975 ;
        RECT 105.530 132.135 110.530 132.305 ;
        RECT 110.820 132.135 115.820 132.305 ;
        RECT 116.110 132.135 121.110 132.305 ;
        RECT 121.400 132.135 126.400 132.305 ;
        RECT 105.300 129.380 105.470 131.920 ;
        RECT 110.590 129.380 110.760 131.920 ;
        RECT 115.880 129.380 116.050 131.920 ;
        RECT 121.170 129.380 121.340 131.920 ;
        RECT 126.460 129.380 126.630 131.920 ;
        RECT 105.530 128.995 110.530 129.165 ;
        RECT 110.820 128.995 115.820 129.165 ;
        RECT 116.110 128.995 121.110 129.165 ;
        RECT 121.400 128.995 126.400 129.165 ;
        RECT 127.625 128.120 128.415 138.400 ;
        RECT 103.705 127.740 128.415 128.120 ;
        RECT 103.705 127.360 130.350 127.740 ;
        RECT 103.775 127.330 130.350 127.360 ;
        RECT 58.830 126.115 72.085 126.250 ;
        RECT 82.775 126.005 95.875 127.285 ;
        RECT 110.465 126.315 121.470 126.925 ;
        RECT 110.465 126.175 121.510 126.315 ;
        RECT 59.310 123.710 101.345 124.645 ;
        RECT 59.310 118.320 60.200 123.710 ;
        RECT 60.970 122.815 70.370 122.985 ;
        RECT 70.660 122.815 80.060 122.985 ;
        RECT 80.350 122.815 89.750 122.985 ;
        RECT 90.040 122.815 99.440 122.985 ;
        RECT 60.740 121.105 60.910 122.645 ;
        RECT 70.430 121.105 70.600 122.645 ;
        RECT 80.120 121.105 80.290 122.645 ;
        RECT 89.810 121.105 89.980 122.645 ;
        RECT 99.500 121.105 99.670 122.645 ;
        RECT 60.970 120.765 70.370 120.935 ;
        RECT 70.660 120.765 80.060 120.935 ;
        RECT 80.350 120.765 89.750 120.935 ;
        RECT 90.040 120.765 99.440 120.935 ;
        RECT 60.740 119.055 60.910 120.595 ;
        RECT 70.430 119.055 70.600 120.595 ;
        RECT 80.120 119.055 80.290 120.595 ;
        RECT 89.810 119.055 89.980 120.595 ;
        RECT 99.500 119.055 99.670 120.595 ;
        RECT 60.970 118.715 70.370 118.885 ;
        RECT 70.660 118.715 80.060 118.885 ;
        RECT 80.350 118.715 89.750 118.885 ;
        RECT 90.040 118.715 99.440 118.885 ;
        RECT 100.500 118.320 101.345 123.710 ;
        RECT 59.310 116.875 101.345 118.320 ;
        RECT 59.355 116.870 101.345 116.875 ;
        RECT 110.500 115.765 110.965 126.175 ;
        RECT 111.455 125.665 113.455 125.835 ;
        RECT 113.745 125.665 115.745 125.835 ;
        RECT 116.035 125.665 118.035 125.835 ;
        RECT 118.325 125.665 120.325 125.835 ;
        RECT 111.225 122.455 111.395 125.495 ;
        RECT 113.515 122.455 113.685 125.495 ;
        RECT 115.805 122.455 115.975 125.495 ;
        RECT 118.095 122.455 118.265 125.495 ;
        RECT 120.385 122.455 120.555 125.495 ;
        RECT 111.455 122.115 113.455 122.285 ;
        RECT 113.745 122.115 115.745 122.285 ;
        RECT 116.035 122.115 118.035 122.285 ;
        RECT 118.325 122.115 120.325 122.285 ;
        RECT 111.455 119.630 113.455 119.800 ;
        RECT 113.745 119.630 115.745 119.800 ;
        RECT 116.035 119.630 118.035 119.800 ;
        RECT 118.325 119.630 120.325 119.800 ;
        RECT 111.225 116.420 111.395 119.460 ;
        RECT 113.515 116.420 113.685 119.460 ;
        RECT 115.805 116.420 115.975 119.460 ;
        RECT 118.095 116.420 118.265 119.460 ;
        RECT 120.385 116.420 120.555 119.460 ;
        RECT 111.455 116.080 113.455 116.250 ;
        RECT 113.745 116.080 115.745 116.250 ;
        RECT 116.035 116.080 118.035 116.250 ;
        RECT 118.325 116.080 120.325 116.250 ;
        RECT 120.900 115.770 121.510 126.175 ;
        RECT 125.930 125.535 130.350 127.330 ;
        RECT 125.930 121.540 126.620 125.535 ;
        RECT 127.195 125.120 127.545 125.290 ;
        RECT 126.965 122.265 127.135 124.905 ;
        RECT 127.605 122.265 127.775 124.905 ;
        RECT 127.195 121.880 127.545 122.050 ;
        RECT 128.175 121.540 128.345 125.535 ;
        RECT 128.975 125.120 129.325 125.290 ;
        RECT 128.745 122.265 128.915 124.905 ;
        RECT 129.385 122.265 129.555 124.905 ;
        RECT 128.975 121.880 129.325 122.050 ;
        RECT 129.935 121.540 130.350 125.535 ;
        RECT 125.930 121.370 130.350 121.540 ;
        RECT 125.930 121.255 126.620 121.370 ;
        RECT 129.935 121.325 130.350 121.370 ;
        RECT 122.940 120.440 130.610 120.830 ;
        RECT 122.940 118.185 126.815 120.440 ;
        RECT 127.305 120.050 127.635 120.220 ;
        RECT 129.085 120.050 129.415 120.220 ;
        RECT 127.165 118.840 127.335 119.880 ;
        RECT 127.605 118.840 127.775 119.880 ;
        RECT 128.945 118.840 129.115 119.880 ;
        RECT 129.385 118.840 129.555 119.880 ;
        RECT 127.305 118.500 127.635 118.670 ;
        RECT 129.085 118.500 129.415 118.670 ;
        RECT 129.880 118.185 130.610 120.440 ;
        RECT 122.940 115.770 130.610 118.185 ;
        RECT 120.900 115.765 130.610 115.770 ;
        RECT 110.270 115.450 130.610 115.765 ;
        RECT 110.270 114.390 123.965 115.450 ;
        RECT 124.445 114.730 126.605 115.080 ;
        RECT 127.645 114.730 129.805 115.080 ;
        RECT 130.255 114.390 130.610 115.450 ;
        RECT 110.270 114.075 130.610 114.390 ;
        RECT 83.360 112.990 86.080 112.995 ;
        RECT 78.540 112.330 82.990 112.945 ;
        RECT 78.540 108.700 79.820 112.330 ;
        RECT 80.400 111.705 81.440 111.875 ;
        RECT 80.060 110.645 80.230 111.645 ;
        RECT 81.610 110.645 81.780 111.645 ;
        RECT 80.400 110.415 81.440 110.585 ;
        RECT 80.060 109.355 80.230 110.355 ;
        RECT 81.610 109.355 81.780 110.355 ;
        RECT 80.400 109.125 81.440 109.295 ;
        RECT 75.775 108.685 79.820 108.700 ;
        RECT 59.875 108.105 79.820 108.685 ;
        RECT 59.875 75.990 61.680 108.105 ;
        RECT 62.310 107.680 66.350 107.850 ;
        RECT 69.715 107.680 73.755 107.850 ;
        RECT 61.970 106.620 62.140 107.620 ;
        RECT 66.520 106.620 66.690 107.620 ;
        RECT 69.375 106.620 69.545 107.620 ;
        RECT 73.925 106.620 74.095 107.620 ;
        RECT 62.310 106.390 66.350 106.560 ;
        RECT 69.715 106.390 73.755 106.560 ;
        RECT 61.970 105.330 62.140 106.330 ;
        RECT 66.520 105.330 66.690 106.330 ;
        RECT 69.375 105.330 69.545 106.330 ;
        RECT 73.925 105.330 74.095 106.330 ;
        RECT 62.310 105.100 66.350 105.270 ;
        RECT 69.715 105.100 73.755 105.270 ;
        RECT 61.970 104.040 62.140 105.040 ;
        RECT 66.520 104.040 66.690 105.040 ;
        RECT 69.375 104.040 69.545 105.040 ;
        RECT 73.925 104.040 74.095 105.040 ;
        RECT 62.310 103.810 66.350 103.980 ;
        RECT 69.715 103.810 73.755 103.980 ;
        RECT 61.970 102.750 62.140 103.750 ;
        RECT 66.520 102.750 66.690 103.750 ;
        RECT 69.375 102.750 69.545 103.750 ;
        RECT 73.925 102.750 74.095 103.750 ;
        RECT 62.310 102.520 66.350 102.690 ;
        RECT 69.715 102.520 73.755 102.690 ;
        RECT 61.970 101.460 62.140 102.460 ;
        RECT 66.520 101.460 66.690 102.460 ;
        RECT 69.375 101.460 69.545 102.460 ;
        RECT 73.925 101.460 74.095 102.460 ;
        RECT 62.310 101.230 66.350 101.400 ;
        RECT 69.715 101.230 73.755 101.400 ;
        RECT 61.970 100.170 62.140 101.170 ;
        RECT 66.520 100.170 66.690 101.170 ;
        RECT 69.375 100.170 69.545 101.170 ;
        RECT 73.925 100.170 74.095 101.170 ;
        RECT 62.310 99.940 66.350 100.110 ;
        RECT 69.715 99.940 73.755 100.110 ;
        RECT 61.970 98.880 62.140 99.880 ;
        RECT 66.520 98.880 66.690 99.880 ;
        RECT 69.375 98.880 69.545 99.880 ;
        RECT 73.925 98.880 74.095 99.880 ;
        RECT 62.310 98.650 66.350 98.820 ;
        RECT 69.715 98.650 73.755 98.820 ;
        RECT 61.970 97.590 62.140 98.590 ;
        RECT 66.520 97.590 66.690 98.590 ;
        RECT 69.375 97.590 69.545 98.590 ;
        RECT 73.925 97.590 74.095 98.590 ;
        RECT 62.310 97.360 66.350 97.530 ;
        RECT 69.715 97.360 73.755 97.530 ;
        RECT 61.970 96.300 62.140 97.300 ;
        RECT 66.520 96.300 66.690 97.300 ;
        RECT 69.375 96.300 69.545 97.300 ;
        RECT 73.925 96.300 74.095 97.300 ;
        RECT 62.310 96.070 66.350 96.240 ;
        RECT 69.715 96.070 73.755 96.240 ;
        RECT 61.970 95.010 62.140 96.010 ;
        RECT 66.520 95.010 66.690 96.010 ;
        RECT 69.375 95.010 69.545 96.010 ;
        RECT 73.925 95.010 74.095 96.010 ;
        RECT 62.310 94.780 66.350 94.950 ;
        RECT 69.715 94.780 73.755 94.950 ;
        RECT 61.970 93.720 62.140 94.720 ;
        RECT 66.520 93.720 66.690 94.720 ;
        RECT 69.375 93.720 69.545 94.720 ;
        RECT 73.925 93.720 74.095 94.720 ;
        RECT 62.310 93.490 66.350 93.660 ;
        RECT 69.715 93.490 73.755 93.660 ;
        RECT 61.970 92.430 62.140 93.430 ;
        RECT 66.520 92.430 66.690 93.430 ;
        RECT 69.375 92.430 69.545 93.430 ;
        RECT 73.925 92.430 74.095 93.430 ;
        RECT 62.310 92.200 66.350 92.370 ;
        RECT 69.715 92.200 73.755 92.370 ;
        RECT 61.970 91.140 62.140 92.140 ;
        RECT 66.520 91.140 66.690 92.140 ;
        RECT 69.375 91.140 69.545 92.140 ;
        RECT 73.925 91.140 74.095 92.140 ;
        RECT 62.310 90.910 66.350 91.080 ;
        RECT 69.715 90.910 73.755 91.080 ;
        RECT 61.970 89.850 62.140 90.850 ;
        RECT 66.520 89.850 66.690 90.850 ;
        RECT 69.375 89.850 69.545 90.850 ;
        RECT 73.925 89.850 74.095 90.850 ;
        RECT 62.310 89.620 66.350 89.790 ;
        RECT 69.715 89.620 73.755 89.790 ;
        RECT 61.970 88.560 62.140 89.560 ;
        RECT 66.520 88.560 66.690 89.560 ;
        RECT 69.375 88.560 69.545 89.560 ;
        RECT 73.925 88.560 74.095 89.560 ;
        RECT 62.310 88.330 66.350 88.500 ;
        RECT 69.715 88.330 73.755 88.500 ;
        RECT 61.970 87.270 62.140 88.270 ;
        RECT 66.520 87.270 66.690 88.270 ;
        RECT 69.375 87.270 69.545 88.270 ;
        RECT 73.925 87.270 74.095 88.270 ;
        RECT 62.310 87.040 66.350 87.210 ;
        RECT 69.715 87.040 73.755 87.210 ;
        RECT 61.970 85.980 62.140 86.980 ;
        RECT 66.520 85.980 66.690 86.980 ;
        RECT 69.375 85.980 69.545 86.980 ;
        RECT 73.925 85.980 74.095 86.980 ;
        RECT 62.310 85.750 66.350 85.920 ;
        RECT 69.715 85.750 73.755 85.920 ;
        RECT 61.970 84.690 62.140 85.690 ;
        RECT 66.520 84.690 66.690 85.690 ;
        RECT 69.375 84.690 69.545 85.690 ;
        RECT 73.925 84.690 74.095 85.690 ;
        RECT 74.710 85.450 79.820 108.105 ;
        RECT 80.060 108.065 80.230 109.065 ;
        RECT 81.610 108.065 81.780 109.065 ;
        RECT 80.400 107.835 81.440 108.005 ;
        RECT 80.060 106.775 80.230 107.775 ;
        RECT 81.610 106.775 81.780 107.775 ;
        RECT 80.400 106.545 81.440 106.715 ;
        RECT 80.060 105.485 80.230 106.485 ;
        RECT 81.610 105.485 81.780 106.485 ;
        RECT 80.400 105.255 81.440 105.425 ;
        RECT 80.060 104.195 80.230 105.195 ;
        RECT 81.610 104.195 81.780 105.195 ;
        RECT 80.400 103.965 81.440 104.135 ;
        RECT 80.060 102.905 80.230 103.905 ;
        RECT 81.610 102.905 81.780 103.905 ;
        RECT 80.400 102.675 81.440 102.845 ;
        RECT 80.060 101.615 80.230 102.615 ;
        RECT 81.610 101.615 81.780 102.615 ;
        RECT 80.400 101.385 81.440 101.555 ;
        RECT 80.060 100.325 80.230 101.325 ;
        RECT 81.610 100.325 81.780 101.325 ;
        RECT 80.400 100.095 81.440 100.265 ;
        RECT 80.060 99.035 80.230 100.035 ;
        RECT 81.610 99.035 81.780 100.035 ;
        RECT 80.400 98.805 81.440 98.975 ;
        RECT 80.060 97.745 80.230 98.745 ;
        RECT 81.610 97.745 81.780 98.745 ;
        RECT 80.400 97.515 81.440 97.685 ;
        RECT 80.060 96.455 80.230 97.455 ;
        RECT 81.610 96.455 81.780 97.455 ;
        RECT 80.400 96.225 81.440 96.395 ;
        RECT 80.060 95.165 80.230 96.165 ;
        RECT 81.610 95.165 81.780 96.165 ;
        RECT 80.400 94.935 81.440 95.105 ;
        RECT 80.060 93.875 80.230 94.875 ;
        RECT 81.610 93.875 81.780 94.875 ;
        RECT 80.400 93.645 81.440 93.815 ;
        RECT 80.060 92.585 80.230 93.585 ;
        RECT 81.610 92.585 81.780 93.585 ;
        RECT 80.400 92.355 81.440 92.525 ;
        RECT 80.060 91.295 80.230 92.295 ;
        RECT 81.610 91.295 81.780 92.295 ;
        RECT 80.400 91.065 81.440 91.235 ;
        RECT 80.060 90.005 80.230 91.005 ;
        RECT 81.610 90.005 81.780 91.005 ;
        RECT 80.400 89.775 81.440 89.945 ;
        RECT 80.060 88.715 80.230 89.715 ;
        RECT 81.610 88.715 81.780 89.715 ;
        RECT 80.400 88.485 81.440 88.655 ;
        RECT 80.060 87.425 80.230 88.425 ;
        RECT 81.610 87.425 81.780 88.425 ;
        RECT 80.400 87.195 81.440 87.365 ;
        RECT 80.060 86.135 80.230 87.135 ;
        RECT 81.610 86.135 81.780 87.135 ;
        RECT 80.400 85.905 81.440 86.075 ;
        RECT 82.295 85.450 82.990 112.330 ;
        RECT 83.360 112.475 88.120 112.990 ;
        RECT 83.360 106.560 83.755 112.475 ;
        RECT 84.335 112.030 85.375 112.200 ;
        RECT 83.950 109.970 84.120 111.970 ;
        RECT 85.590 109.970 85.760 111.970 ;
        RECT 84.335 109.740 85.375 109.910 ;
        RECT 84.335 109.125 85.375 109.295 ;
        RECT 83.950 107.065 84.120 109.065 ;
        RECT 85.590 107.065 85.760 109.065 ;
        RECT 84.335 106.835 85.375 107.005 ;
        RECT 86.000 106.560 88.120 112.475 ;
        RECT 110.285 109.725 112.700 114.075 ;
        RECT 113.250 113.580 118.790 113.750 ;
        RECT 112.910 112.020 113.080 113.520 ;
        RECT 118.960 112.020 119.130 113.520 ;
        RECT 113.250 111.790 118.790 111.960 ;
        RECT 112.910 110.230 113.080 111.730 ;
        RECT 118.960 110.230 119.130 111.730 ;
        RECT 113.250 110.000 118.790 110.170 ;
        RECT 119.470 109.725 121.050 114.075 ;
        RECT 121.415 114.070 130.610 114.075 ;
        RECT 110.285 107.825 121.050 109.725 ;
        RECT 83.360 106.145 88.120 106.560 ;
        RECT 83.370 106.135 88.120 106.145 ;
        RECT 84.190 103.595 88.120 106.135 ;
        RECT 83.315 103.115 88.120 103.595 ;
        RECT 83.315 100.130 83.730 103.115 ;
        RECT 85.995 103.110 88.120 103.115 ;
        RECT 84.335 102.675 85.375 102.845 ;
        RECT 83.950 100.615 84.120 102.615 ;
        RECT 85.590 100.615 85.760 102.615 ;
        RECT 86.000 100.610 88.120 103.110 ;
        RECT 84.335 100.385 85.375 100.555 ;
        RECT 85.995 100.130 88.120 100.610 ;
        RECT 83.315 99.675 88.120 100.130 ;
        RECT 84.190 97.145 88.120 99.675 ;
        RECT 83.360 96.745 88.120 97.145 ;
        RECT 83.360 93.640 83.740 96.745 ;
        RECT 84.335 96.225 85.375 96.395 ;
        RECT 83.950 94.165 84.120 96.165 ;
        RECT 85.590 94.165 85.760 96.165 ;
        RECT 84.335 93.935 85.375 94.105 ;
        RECT 86.000 93.640 88.120 96.745 ;
        RECT 83.360 93.215 88.120 93.640 ;
        RECT 83.360 93.195 83.740 93.215 ;
        RECT 83.330 90.640 83.670 90.645 ;
        RECT 84.250 90.640 88.120 93.215 ;
        RECT 83.330 90.250 88.120 90.640 ;
        RECT 83.330 87.190 83.670 90.250 ;
        RECT 84.335 89.775 85.375 89.945 ;
        RECT 83.950 87.715 84.120 89.715 ;
        RECT 85.590 87.715 85.760 89.715 ;
        RECT 84.335 87.485 85.375 87.655 ;
        RECT 86.000 87.190 88.120 90.250 ;
        RECT 83.330 86.810 88.120 87.190 ;
        RECT 83.340 86.800 88.120 86.810 ;
        RECT 74.710 84.835 82.990 85.450 ;
        RECT 85.960 85.085 88.120 86.800 ;
        RECT 83.485 84.840 88.120 85.085 ;
        RECT 74.710 84.810 78.595 84.835 ;
        RECT 62.310 84.460 66.350 84.630 ;
        RECT 69.715 84.460 73.755 84.630 ;
        RECT 61.970 83.400 62.140 84.400 ;
        RECT 66.520 83.400 66.690 84.400 ;
        RECT 69.375 83.400 69.545 84.400 ;
        RECT 73.925 83.400 74.095 84.400 ;
        RECT 62.310 83.170 66.350 83.340 ;
        RECT 69.715 83.170 73.755 83.340 ;
        RECT 61.970 82.110 62.140 83.110 ;
        RECT 66.520 82.110 66.690 83.110 ;
        RECT 69.375 82.110 69.545 83.110 ;
        RECT 73.925 82.110 74.095 83.110 ;
        RECT 62.310 81.880 66.350 82.050 ;
        RECT 69.715 81.880 73.755 82.050 ;
        RECT 74.710 81.960 76.210 84.810 ;
        RECT 61.970 80.820 62.140 81.820 ;
        RECT 66.520 80.820 66.690 81.820 ;
        RECT 69.375 80.820 69.545 81.820 ;
        RECT 73.925 80.820 74.095 81.820 ;
        RECT 74.710 80.785 82.620 81.960 ;
        RECT 62.310 80.590 66.350 80.760 ;
        RECT 69.715 80.590 73.755 80.760 ;
        RECT 61.970 79.530 62.140 80.530 ;
        RECT 66.520 79.530 66.690 80.530 ;
        RECT 69.375 79.530 69.545 80.530 ;
        RECT 73.925 79.530 74.095 80.530 ;
        RECT 62.310 79.300 66.350 79.470 ;
        RECT 69.715 79.300 73.755 79.470 ;
        RECT 61.970 78.240 62.140 79.240 ;
        RECT 66.520 78.240 66.690 79.240 ;
        RECT 69.375 78.240 69.545 79.240 ;
        RECT 73.925 78.240 74.095 79.240 ;
        RECT 62.310 78.010 66.350 78.180 ;
        RECT 69.715 78.010 73.755 78.180 ;
        RECT 61.970 76.950 62.140 77.950 ;
        RECT 66.520 76.950 66.690 77.950 ;
        RECT 69.375 76.950 69.545 77.950 ;
        RECT 73.925 76.950 74.095 77.950 ;
        RECT 62.310 76.720 66.350 76.890 ;
        RECT 69.715 76.720 73.755 76.890 ;
        RECT 74.710 76.790 77.355 80.785 ;
        RECT 77.665 77.005 81.135 80.475 ;
        RECT 74.745 76.695 77.355 76.790 ;
        RECT 81.445 76.695 82.620 80.785 ;
        RECT 74.745 75.990 82.620 76.695 ;
        RECT 59.875 75.530 82.620 75.990 ;
        RECT 59.875 75.095 61.680 75.530 ;
        RECT 75.750 75.525 82.620 75.530 ;
        RECT 76.180 75.520 82.620 75.525 ;
        RECT 83.485 75.640 83.725 84.840 ;
        RECT 85.960 84.625 88.120 84.840 ;
        RECT 84.335 84.335 85.375 84.505 ;
        RECT 83.950 83.275 84.120 84.275 ;
        RECT 85.590 83.275 85.760 84.275 ;
        RECT 84.335 83.045 85.375 83.215 ;
        RECT 83.950 81.985 84.120 82.985 ;
        RECT 85.590 81.985 85.760 82.985 ;
        RECT 84.335 81.755 85.375 81.925 ;
        RECT 85.960 81.365 88.115 84.625 ;
        RECT 84.335 80.710 84.875 80.880 ;
        RECT 83.950 78.650 84.120 80.650 ;
        RECT 85.090 78.650 85.260 80.650 ;
        RECT 84.335 78.420 84.875 78.590 ;
        RECT 83.950 76.360 84.120 78.360 ;
        RECT 85.090 76.360 85.260 78.360 ;
        RECT 85.945 76.425 88.115 81.365 ;
        RECT 84.335 76.130 84.875 76.300 ;
        RECT 85.950 76.195 88.115 76.425 ;
        RECT 85.945 75.640 88.115 76.195 ;
        RECT 83.485 75.380 88.115 75.640 ;
        RECT 85.945 74.995 88.115 75.380 ;
        RECT 88.630 54.010 129.510 55.700 ;
        RECT 13.050 52.115 14.855 52.550 ;
        RECT 39.120 52.265 41.290 52.650 ;
        RECT 29.355 52.120 35.795 52.125 ;
        RECT 28.925 52.115 35.795 52.120 ;
        RECT 13.050 51.655 35.795 52.115 ;
        RECT 13.050 19.540 14.855 51.655 ;
        RECT 27.920 50.950 35.795 51.655 ;
        RECT 15.485 50.755 19.525 50.925 ;
        RECT 22.890 50.755 26.930 50.925 ;
        RECT 27.920 50.855 30.530 50.950 ;
        RECT 15.145 49.695 15.315 50.695 ;
        RECT 19.695 49.695 19.865 50.695 ;
        RECT 22.550 49.695 22.720 50.695 ;
        RECT 27.100 49.695 27.270 50.695 ;
        RECT 15.485 49.465 19.525 49.635 ;
        RECT 22.890 49.465 26.930 49.635 ;
        RECT 15.145 48.405 15.315 49.405 ;
        RECT 19.695 48.405 19.865 49.405 ;
        RECT 22.550 48.405 22.720 49.405 ;
        RECT 27.100 48.405 27.270 49.405 ;
        RECT 15.485 48.175 19.525 48.345 ;
        RECT 22.890 48.175 26.930 48.345 ;
        RECT 15.145 47.115 15.315 48.115 ;
        RECT 19.695 47.115 19.865 48.115 ;
        RECT 22.550 47.115 22.720 48.115 ;
        RECT 27.100 47.115 27.270 48.115 ;
        RECT 15.485 46.885 19.525 47.055 ;
        RECT 22.890 46.885 26.930 47.055 ;
        RECT 27.885 46.860 30.530 50.855 ;
        RECT 30.840 47.170 34.310 50.640 ;
        RECT 34.620 46.860 35.795 50.950 ;
        RECT 15.145 45.825 15.315 46.825 ;
        RECT 19.695 45.825 19.865 46.825 ;
        RECT 22.550 45.825 22.720 46.825 ;
        RECT 27.100 45.825 27.270 46.825 ;
        RECT 15.485 45.595 19.525 45.765 ;
        RECT 22.890 45.595 26.930 45.765 ;
        RECT 27.885 45.685 35.795 46.860 ;
        RECT 36.660 52.005 41.290 52.265 ;
        RECT 15.145 44.535 15.315 45.535 ;
        RECT 19.695 44.535 19.865 45.535 ;
        RECT 22.550 44.535 22.720 45.535 ;
        RECT 27.100 44.535 27.270 45.535 ;
        RECT 15.485 44.305 19.525 44.475 ;
        RECT 22.890 44.305 26.930 44.475 ;
        RECT 15.145 43.245 15.315 44.245 ;
        RECT 19.695 43.245 19.865 44.245 ;
        RECT 22.550 43.245 22.720 44.245 ;
        RECT 27.100 43.245 27.270 44.245 ;
        RECT 15.485 43.015 19.525 43.185 ;
        RECT 22.890 43.015 26.930 43.185 ;
        RECT 15.145 41.955 15.315 42.955 ;
        RECT 19.695 41.955 19.865 42.955 ;
        RECT 22.550 41.955 22.720 42.955 ;
        RECT 27.100 41.955 27.270 42.955 ;
        RECT 27.885 42.320 29.385 45.685 ;
        RECT 36.660 42.805 36.900 52.005 ;
        RECT 37.510 51.345 38.050 51.515 ;
        RECT 39.120 51.450 41.290 52.005 ;
        RECT 37.125 49.285 37.295 51.285 ;
        RECT 38.265 49.285 38.435 51.285 ;
        RECT 39.125 51.220 41.290 51.450 ;
        RECT 37.510 49.055 38.050 49.225 ;
        RECT 37.125 46.995 37.295 48.995 ;
        RECT 38.265 46.995 38.435 48.995 ;
        RECT 37.510 46.765 38.050 46.935 ;
        RECT 39.120 46.280 41.290 51.220 ;
        RECT 88.630 48.165 89.900 54.010 ;
        RECT 91.105 53.565 109.105 53.735 ;
        RECT 109.395 53.565 127.395 53.735 ;
        RECT 90.875 51.510 91.045 53.350 ;
        RECT 109.165 51.510 109.335 53.350 ;
        RECT 127.455 51.510 127.625 53.350 ;
        RECT 91.105 51.125 109.105 51.295 ;
        RECT 109.395 51.125 127.395 51.295 ;
        RECT 90.875 49.070 91.045 50.910 ;
        RECT 109.165 49.070 109.335 50.910 ;
        RECT 127.455 49.070 127.625 50.910 ;
        RECT 91.105 48.685 109.105 48.855 ;
        RECT 109.395 48.685 127.395 48.855 ;
        RECT 128.460 48.165 129.505 54.010 ;
        RECT 88.630 47.500 129.505 48.165 ;
        RECT 37.510 45.720 38.550 45.890 ;
        RECT 37.125 44.660 37.295 45.660 ;
        RECT 38.765 44.660 38.935 45.660 ;
        RECT 37.510 44.430 38.550 44.600 ;
        RECT 37.125 43.370 37.295 44.370 ;
        RECT 38.765 43.370 38.935 44.370 ;
        RECT 37.510 43.140 38.550 43.310 ;
        RECT 39.135 42.805 41.290 46.280 ;
        RECT 36.660 42.560 41.290 42.805 ;
        RECT 39.135 42.385 41.290 42.560 ;
        RECT 88.635 44.625 124.380 45.325 ;
        RECT 27.885 42.315 31.760 42.320 ;
        RECT 15.485 41.725 19.525 41.895 ;
        RECT 22.890 41.725 26.930 41.895 ;
        RECT 27.885 41.700 36.165 42.315 ;
        RECT 15.145 40.665 15.315 41.665 ;
        RECT 19.695 40.665 19.865 41.665 ;
        RECT 22.550 40.665 22.720 41.665 ;
        RECT 27.100 40.665 27.270 41.665 ;
        RECT 15.485 40.435 19.525 40.605 ;
        RECT 22.890 40.435 26.930 40.605 ;
        RECT 15.145 39.375 15.315 40.375 ;
        RECT 19.695 39.375 19.865 40.375 ;
        RECT 22.550 39.375 22.720 40.375 ;
        RECT 27.100 39.375 27.270 40.375 ;
        RECT 15.485 39.145 19.525 39.315 ;
        RECT 22.890 39.145 26.930 39.315 ;
        RECT 15.145 38.085 15.315 39.085 ;
        RECT 19.695 38.085 19.865 39.085 ;
        RECT 22.550 38.085 22.720 39.085 ;
        RECT 27.100 38.085 27.270 39.085 ;
        RECT 15.485 37.855 19.525 38.025 ;
        RECT 22.890 37.855 26.930 38.025 ;
        RECT 15.145 36.795 15.315 37.795 ;
        RECT 19.695 36.795 19.865 37.795 ;
        RECT 22.550 36.795 22.720 37.795 ;
        RECT 27.100 36.795 27.270 37.795 ;
        RECT 15.485 36.565 19.525 36.735 ;
        RECT 22.890 36.565 26.930 36.735 ;
        RECT 15.145 35.505 15.315 36.505 ;
        RECT 19.695 35.505 19.865 36.505 ;
        RECT 22.550 35.505 22.720 36.505 ;
        RECT 27.100 35.505 27.270 36.505 ;
        RECT 15.485 35.275 19.525 35.445 ;
        RECT 22.890 35.275 26.930 35.445 ;
        RECT 15.145 34.215 15.315 35.215 ;
        RECT 19.695 34.215 19.865 35.215 ;
        RECT 22.550 34.215 22.720 35.215 ;
        RECT 27.100 34.215 27.270 35.215 ;
        RECT 15.485 33.985 19.525 34.155 ;
        RECT 22.890 33.985 26.930 34.155 ;
        RECT 15.145 32.925 15.315 33.925 ;
        RECT 19.695 32.925 19.865 33.925 ;
        RECT 22.550 32.925 22.720 33.925 ;
        RECT 27.100 32.925 27.270 33.925 ;
        RECT 15.485 32.695 19.525 32.865 ;
        RECT 22.890 32.695 26.930 32.865 ;
        RECT 15.145 31.635 15.315 32.635 ;
        RECT 19.695 31.635 19.865 32.635 ;
        RECT 22.550 31.635 22.720 32.635 ;
        RECT 27.100 31.635 27.270 32.635 ;
        RECT 15.485 31.405 19.525 31.575 ;
        RECT 22.890 31.405 26.930 31.575 ;
        RECT 15.145 30.345 15.315 31.345 ;
        RECT 19.695 30.345 19.865 31.345 ;
        RECT 22.550 30.345 22.720 31.345 ;
        RECT 27.100 30.345 27.270 31.345 ;
        RECT 15.485 30.115 19.525 30.285 ;
        RECT 22.890 30.115 26.930 30.285 ;
        RECT 15.145 29.055 15.315 30.055 ;
        RECT 19.695 29.055 19.865 30.055 ;
        RECT 22.550 29.055 22.720 30.055 ;
        RECT 27.100 29.055 27.270 30.055 ;
        RECT 15.485 28.825 19.525 28.995 ;
        RECT 22.890 28.825 26.930 28.995 ;
        RECT 15.145 27.765 15.315 28.765 ;
        RECT 19.695 27.765 19.865 28.765 ;
        RECT 22.550 27.765 22.720 28.765 ;
        RECT 27.100 27.765 27.270 28.765 ;
        RECT 15.485 27.535 19.525 27.705 ;
        RECT 22.890 27.535 26.930 27.705 ;
        RECT 15.145 26.475 15.315 27.475 ;
        RECT 19.695 26.475 19.865 27.475 ;
        RECT 22.550 26.475 22.720 27.475 ;
        RECT 27.100 26.475 27.270 27.475 ;
        RECT 15.485 26.245 19.525 26.415 ;
        RECT 22.890 26.245 26.930 26.415 ;
        RECT 15.145 25.185 15.315 26.185 ;
        RECT 19.695 25.185 19.865 26.185 ;
        RECT 22.550 25.185 22.720 26.185 ;
        RECT 27.100 25.185 27.270 26.185 ;
        RECT 15.485 24.955 19.525 25.125 ;
        RECT 22.890 24.955 26.930 25.125 ;
        RECT 15.145 23.895 15.315 24.895 ;
        RECT 19.695 23.895 19.865 24.895 ;
        RECT 22.550 23.895 22.720 24.895 ;
        RECT 27.100 23.895 27.270 24.895 ;
        RECT 15.485 23.665 19.525 23.835 ;
        RECT 22.890 23.665 26.930 23.835 ;
        RECT 15.145 22.605 15.315 23.605 ;
        RECT 19.695 22.605 19.865 23.605 ;
        RECT 22.550 22.605 22.720 23.605 ;
        RECT 27.100 22.605 27.270 23.605 ;
        RECT 15.485 22.375 19.525 22.545 ;
        RECT 22.890 22.375 26.930 22.545 ;
        RECT 15.145 21.315 15.315 22.315 ;
        RECT 19.695 21.315 19.865 22.315 ;
        RECT 22.550 21.315 22.720 22.315 ;
        RECT 27.100 21.315 27.270 22.315 ;
        RECT 15.485 21.085 19.525 21.255 ;
        RECT 22.890 21.085 26.930 21.255 ;
        RECT 15.145 20.025 15.315 21.025 ;
        RECT 19.695 20.025 19.865 21.025 ;
        RECT 22.550 20.025 22.720 21.025 ;
        RECT 27.100 20.025 27.270 21.025 ;
        RECT 15.485 19.795 19.525 19.965 ;
        RECT 22.890 19.795 26.930 19.965 ;
        RECT 27.885 19.540 32.995 41.700 ;
        RECT 33.575 41.075 34.615 41.245 ;
        RECT 33.235 40.015 33.405 41.015 ;
        RECT 34.785 40.015 34.955 41.015 ;
        RECT 33.575 39.785 34.615 39.955 ;
        RECT 33.235 38.725 33.405 39.725 ;
        RECT 34.785 38.725 34.955 39.725 ;
        RECT 33.575 38.495 34.615 38.665 ;
        RECT 33.235 37.435 33.405 38.435 ;
        RECT 34.785 37.435 34.955 38.435 ;
        RECT 33.575 37.205 34.615 37.375 ;
        RECT 33.235 36.145 33.405 37.145 ;
        RECT 34.785 36.145 34.955 37.145 ;
        RECT 33.575 35.915 34.615 36.085 ;
        RECT 33.235 34.855 33.405 35.855 ;
        RECT 34.785 34.855 34.955 35.855 ;
        RECT 33.575 34.625 34.615 34.795 ;
        RECT 33.235 33.565 33.405 34.565 ;
        RECT 34.785 33.565 34.955 34.565 ;
        RECT 33.575 33.335 34.615 33.505 ;
        RECT 33.235 32.275 33.405 33.275 ;
        RECT 34.785 32.275 34.955 33.275 ;
        RECT 33.575 32.045 34.615 32.215 ;
        RECT 33.235 30.985 33.405 31.985 ;
        RECT 34.785 30.985 34.955 31.985 ;
        RECT 33.575 30.755 34.615 30.925 ;
        RECT 33.235 29.695 33.405 30.695 ;
        RECT 34.785 29.695 34.955 30.695 ;
        RECT 33.575 29.465 34.615 29.635 ;
        RECT 33.235 28.405 33.405 29.405 ;
        RECT 34.785 28.405 34.955 29.405 ;
        RECT 33.575 28.175 34.615 28.345 ;
        RECT 33.235 27.115 33.405 28.115 ;
        RECT 34.785 27.115 34.955 28.115 ;
        RECT 33.575 26.885 34.615 27.055 ;
        RECT 33.235 25.825 33.405 26.825 ;
        RECT 34.785 25.825 34.955 26.825 ;
        RECT 33.575 25.595 34.615 25.765 ;
        RECT 33.235 24.535 33.405 25.535 ;
        RECT 34.785 24.535 34.955 25.535 ;
        RECT 33.575 24.305 34.615 24.475 ;
        RECT 33.235 23.245 33.405 24.245 ;
        RECT 34.785 23.245 34.955 24.245 ;
        RECT 33.575 23.015 34.615 23.185 ;
        RECT 33.235 21.955 33.405 22.955 ;
        RECT 34.785 21.955 34.955 22.955 ;
        RECT 33.575 21.725 34.615 21.895 ;
        RECT 33.235 20.665 33.405 21.665 ;
        RECT 34.785 20.665 34.955 21.665 ;
        RECT 33.575 20.435 34.615 20.605 ;
        RECT 13.050 18.960 32.995 19.540 ;
        RECT 33.235 19.375 33.405 20.375 ;
        RECT 34.785 19.375 34.955 20.375 ;
        RECT 33.575 19.145 34.615 19.315 ;
        RECT 31.715 14.820 32.995 18.960 ;
        RECT 33.235 18.085 33.405 19.085 ;
        RECT 34.785 18.085 34.955 19.085 ;
        RECT 33.575 17.855 34.615 18.025 ;
        RECT 33.235 16.795 33.405 17.795 ;
        RECT 34.785 16.795 34.955 17.795 ;
        RECT 33.575 16.565 34.615 16.735 ;
        RECT 33.235 15.505 33.405 16.505 ;
        RECT 34.785 15.505 34.955 16.505 ;
        RECT 33.575 15.275 34.615 15.445 ;
        RECT 35.470 14.820 36.165 41.700 ;
        RECT 36.515 40.340 40.800 40.350 ;
        RECT 36.505 39.960 40.800 40.340 ;
        RECT 36.505 36.900 36.845 39.960 ;
        RECT 37.510 39.495 38.550 39.665 ;
        RECT 37.125 37.435 37.295 39.435 ;
        RECT 38.765 37.435 38.935 39.435 ;
        RECT 37.510 37.205 38.550 37.375 ;
        RECT 39.175 36.900 40.800 39.960 ;
        RECT 88.635 36.920 96.015 44.625 ;
        RECT 97.155 44.160 109.155 44.330 ;
        RECT 109.445 44.160 121.445 44.330 ;
        RECT 96.925 37.950 97.095 43.990 ;
        RECT 109.215 37.950 109.385 43.990 ;
        RECT 121.505 37.950 121.675 43.990 ;
        RECT 97.155 37.610 109.155 37.780 ;
        RECT 109.445 37.610 121.445 37.780 ;
        RECT 36.505 36.510 40.800 36.900 ;
        RECT 36.505 36.505 36.845 36.510 ;
        RECT 36.535 33.935 36.915 33.955 ;
        RECT 37.425 33.935 40.800 36.510 ;
        RECT 36.535 33.510 40.800 33.935 ;
        RECT 36.535 30.405 36.915 33.510 ;
        RECT 37.510 33.045 38.550 33.215 ;
        RECT 37.125 30.985 37.295 32.985 ;
        RECT 38.765 30.985 38.935 32.985 ;
        RECT 37.510 30.755 38.550 30.925 ;
        RECT 39.175 30.405 40.800 33.510 ;
        RECT 36.535 30.005 40.800 30.405 ;
        RECT 37.365 27.475 40.800 30.005 ;
        RECT 88.630 36.735 96.015 36.920 ;
        RECT 88.630 30.505 89.685 36.735 ;
        RECT 90.210 36.175 93.250 36.345 ;
        RECT 89.870 31.115 90.040 36.115 ;
        RECT 93.420 31.115 93.590 36.115 ;
        RECT 90.210 30.505 93.250 31.055 ;
        RECT 93.890 30.505 96.015 36.735 ;
        RECT 97.150 34.785 109.150 34.955 ;
        RECT 109.440 34.785 121.440 34.955 ;
        RECT 88.630 29.355 96.015 30.505 ;
        RECT 36.490 27.020 40.800 27.475 ;
        RECT 36.490 24.035 36.905 27.020 ;
        RECT 37.510 26.595 38.550 26.765 ;
        RECT 39.170 26.540 40.800 27.020 ;
        RECT 37.125 24.535 37.295 26.535 ;
        RECT 38.765 24.535 38.935 26.535 ;
        RECT 37.510 24.305 38.550 24.475 ;
        RECT 39.175 24.040 40.800 26.540 ;
        RECT 88.620 27.955 96.015 29.355 ;
        RECT 96.920 28.575 97.090 34.615 ;
        RECT 109.210 28.575 109.380 34.615 ;
        RECT 121.500 28.575 121.670 34.615 ;
        RECT 97.150 28.235 109.150 28.405 ;
        RECT 109.440 28.235 121.440 28.405 ;
        RECT 122.630 27.955 124.380 44.625 ;
        RECT 88.620 26.405 124.380 27.955 ;
        RECT 39.170 24.035 40.800 24.040 ;
        RECT 36.490 23.555 40.800 24.035 ;
        RECT 37.365 21.370 40.800 23.555 ;
        RECT 37.365 21.015 40.805 21.370 ;
        RECT 36.545 21.005 40.805 21.015 ;
        RECT 31.715 14.205 36.165 14.820 ;
        RECT 36.535 20.590 40.805 21.005 ;
        RECT 36.535 14.675 36.930 20.590 ;
        RECT 37.510 20.145 38.550 20.315 ;
        RECT 37.125 18.085 37.295 20.085 ;
        RECT 38.765 18.085 38.935 20.085 ;
        RECT 37.510 17.855 38.550 18.025 ;
        RECT 37.510 17.240 38.550 17.410 ;
        RECT 37.125 15.180 37.295 17.180 ;
        RECT 38.765 15.180 38.935 17.180 ;
        RECT 37.510 14.950 38.550 15.120 ;
        RECT 39.175 14.675 40.805 20.590 ;
        RECT 36.535 14.160 40.805 14.675 ;
        RECT 36.535 14.155 39.255 14.160 ;
      LAYER met1 ;
        RECT 58.940 164.015 72.020 165.090 ;
        RECT 16.945 153.975 56.055 154.480 ;
        RECT 17.595 152.465 54.830 152.695 ;
        RECT 17.595 150.455 18.595 152.465 ;
        RECT 17.595 145.300 18.025 150.455 ;
        RECT 19.480 150.255 35.675 152.465 ;
        RECT 36.590 152.200 36.820 152.260 ;
        RECT 36.520 150.520 36.890 152.200 ;
        RECT 36.590 150.460 36.820 150.520 ;
        RECT 37.790 150.255 53.985 152.465 ;
        RECT 54.810 150.465 55.820 152.265 ;
        RECT 54.880 150.460 55.110 150.465 ;
        RECT 18.580 150.025 36.540 150.255 ;
        RECT 36.870 150.025 54.830 150.255 ;
        RECT 18.165 148.015 18.595 149.820 ;
        RECT 19.480 147.815 35.675 150.025 ;
        RECT 36.590 149.760 36.820 149.820 ;
        RECT 36.520 148.080 36.890 149.760 ;
        RECT 36.590 148.020 36.820 148.080 ;
        RECT 37.790 147.815 53.985 150.025 ;
        RECT 54.820 147.815 55.250 149.820 ;
        RECT 18.580 147.585 55.250 147.815 ;
        RECT 55.390 146.225 55.820 150.465 ;
        RECT 58.950 147.005 59.875 164.015 ;
        RECT 60.940 162.845 62.800 163.075 ;
        RECT 63.130 162.845 64.990 163.075 ;
        RECT 65.320 162.845 67.180 163.075 ;
        RECT 67.510 162.845 69.370 163.075 ;
        RECT 60.660 152.700 60.890 162.640 ;
        RECT 60.560 147.700 60.980 152.700 ;
        RECT 60.660 147.640 60.890 147.700 ;
        RECT 61.300 147.450 62.325 162.845 ;
        RECT 62.850 162.580 63.080 162.640 ;
        RECT 62.735 159.580 63.195 162.580 ;
        RECT 62.850 147.640 63.080 159.580 ;
        RECT 63.565 147.450 64.590 162.845 ;
        RECT 65.040 158.885 65.270 162.640 ;
        RECT 64.945 153.885 65.365 158.885 ;
        RECT 65.040 147.640 65.270 153.885 ;
        RECT 65.745 147.450 66.770 162.845 ;
        RECT 67.230 162.580 67.460 162.640 ;
        RECT 67.115 159.580 67.575 162.580 ;
        RECT 67.230 147.640 67.460 159.580 ;
        RECT 67.945 147.450 68.970 162.845 ;
        RECT 69.420 152.700 69.650 162.640 ;
        RECT 69.325 147.700 69.745 152.700 ;
        RECT 70.870 148.690 71.640 161.210 ;
        RECT 69.420 147.640 69.650 147.700 ;
        RECT 60.950 147.435 62.450 147.450 ;
        RECT 63.140 147.435 64.640 147.450 ;
        RECT 65.330 147.435 66.830 147.450 ;
        RECT 67.520 147.435 69.020 147.450 ;
        RECT 60.940 147.205 62.800 147.435 ;
        RECT 63.130 147.205 64.990 147.435 ;
        RECT 65.320 147.205 67.180 147.435 ;
        RECT 67.510 147.205 69.370 147.435 ;
        RECT 60.950 147.190 62.450 147.205 ;
        RECT 63.140 147.190 64.640 147.205 ;
        RECT 65.330 147.190 66.830 147.205 ;
        RECT 67.520 147.190 69.020 147.205 ;
        RECT 58.970 146.945 59.855 147.005 ;
        RECT 18.165 145.725 78.155 146.225 ;
        RECT 17.595 144.800 55.300 145.300 ;
        RECT 54.870 144.680 55.300 144.800 ;
        RECT 54.870 144.180 70.095 144.680 ;
        RECT 24.630 143.060 36.590 143.290 ;
        RECT 36.920 143.060 48.880 143.290 ;
        RECT 61.290 143.190 62.790 143.205 ;
        RECT 63.480 143.190 64.980 143.205 ;
        RECT 65.670 143.190 67.170 143.205 ;
        RECT 67.860 143.190 69.360 143.205 ;
        RECT 24.350 142.840 24.580 142.900 ;
        RECT 24.110 137.170 24.640 142.840 ;
        RECT 24.350 136.900 24.580 137.170 ;
        RECT 27.870 136.770 33.295 143.060 ;
        RECT 36.640 138.715 36.870 142.900 ;
        RECT 36.580 137.120 36.940 138.715 ;
        RECT 36.640 136.900 36.870 137.120 ;
        RECT 40.390 136.770 45.825 143.060 ;
        RECT 59.055 142.915 59.855 142.975 ;
        RECT 60.940 142.960 62.800 143.190 ;
        RECT 63.130 142.960 64.990 143.190 ;
        RECT 65.320 142.960 67.180 143.190 ;
        RECT 67.510 142.960 69.370 143.190 ;
        RECT 61.290 142.945 62.790 142.960 ;
        RECT 63.480 142.945 64.980 142.960 ;
        RECT 65.670 142.945 67.170 142.960 ;
        RECT 67.860 142.945 69.360 142.960 ;
        RECT 48.930 142.840 49.160 142.900 ;
        RECT 48.870 137.235 49.400 142.840 ;
        RECT 48.930 136.900 49.160 137.235 ;
        RECT 24.660 136.740 36.580 136.770 ;
        RECT 36.930 136.740 48.870 136.770 ;
        RECT 24.630 136.510 36.590 136.740 ;
        RECT 36.920 136.510 48.880 136.740 ;
        RECT 24.660 136.485 36.580 136.510 ;
        RECT 36.930 136.485 48.870 136.510 ;
        RECT 24.710 135.805 38.025 136.200 ;
        RECT 17.695 135.305 20.675 135.360 ;
        RECT 17.685 135.075 20.685 135.305 ;
        RECT 17.295 134.030 17.525 135.025 ;
        RECT 20.845 134.120 21.140 135.025 ;
        RECT 35.475 134.270 48.820 134.715 ;
        RECT 20.785 134.030 21.145 134.120 ;
        RECT 17.295 131.045 21.145 134.030 ;
        RECT 24.635 133.915 36.575 133.945 ;
        RECT 36.925 133.915 48.865 133.940 ;
        RECT 24.625 133.685 36.585 133.915 ;
        RECT 36.915 133.685 48.875 133.915 ;
        RECT 24.635 133.660 36.575 133.685 ;
        RECT 24.345 133.465 24.575 133.525 ;
        RECT 17.295 130.065 17.525 131.045 ;
        RECT 20.785 130.125 21.145 131.045 ;
        RECT 20.845 130.065 21.140 130.125 ;
        RECT 17.685 129.785 20.685 130.015 ;
        RECT 23.580 127.760 24.635 133.465 ;
        RECT 24.345 127.525 24.575 127.760 ;
        RECT 27.845 127.370 33.280 133.660 ;
        RECT 36.925 133.655 48.865 133.685 ;
        RECT 36.635 133.310 36.865 133.525 ;
        RECT 36.575 131.715 36.935 133.310 ;
        RECT 36.635 127.525 36.865 131.715 ;
        RECT 16.555 126.765 19.440 127.295 ;
        RECT 24.625 127.110 36.585 127.370 ;
        RECT 36.925 127.365 39.425 127.375 ;
        RECT 40.345 127.365 45.780 133.655 ;
        RECT 48.925 133.465 49.155 133.525 ;
        RECT 48.860 128.105 49.720 133.465 ;
        RECT 48.925 127.525 49.155 128.105 ;
        RECT 36.915 127.135 48.875 127.365 ;
        RECT 36.925 127.115 39.425 127.135 ;
        RECT 59.035 127.035 59.875 142.915 ;
        RECT 60.660 142.695 60.890 142.755 ;
        RECT 60.565 137.695 60.985 142.695 ;
        RECT 60.660 127.755 60.890 137.695 ;
        RECT 61.320 127.550 62.345 142.945 ;
        RECT 62.850 130.815 63.080 142.755 ;
        RECT 62.735 127.815 63.195 130.815 ;
        RECT 62.850 127.755 63.080 127.815 ;
        RECT 63.585 127.550 64.610 142.945 ;
        RECT 65.040 136.895 65.270 142.755 ;
        RECT 64.945 131.895 65.365 136.895 ;
        RECT 65.040 127.755 65.270 131.895 ;
        RECT 65.765 127.550 66.790 142.945 ;
        RECT 67.230 130.815 67.460 142.755 ;
        RECT 67.110 127.815 67.570 130.815 ;
        RECT 67.230 127.755 67.460 127.815 ;
        RECT 67.925 127.550 68.950 142.945 ;
        RECT 69.420 142.695 69.650 142.755 ;
        RECT 69.325 137.695 69.745 142.695 ;
        RECT 126.985 140.815 128.340 140.850 ;
        RECT 103.440 140.790 128.340 140.815 ;
        RECT 69.420 127.755 69.650 137.695 ;
        RECT 70.950 137.525 71.720 140.045 ;
        RECT 103.440 138.965 128.360 140.790 ;
        RECT 103.440 138.930 128.340 138.965 ;
        RECT 94.225 137.525 95.720 137.550 ;
        RECT 70.950 137.490 95.720 137.525 ;
        RECT 70.950 136.005 95.740 137.490 ;
        RECT 60.940 127.320 62.800 127.550 ;
        RECT 63.130 127.320 64.990 127.550 ;
        RECT 65.320 127.320 67.180 127.550 ;
        RECT 67.510 127.320 69.370 127.550 ;
        RECT 70.950 127.525 71.720 136.005 ;
        RECT 59.030 126.900 59.875 127.035 ;
        RECT 82.970 127.285 84.195 136.005 ;
        RECT 85.085 135.190 86.845 135.420 ;
        RECT 87.175 135.190 88.935 135.420 ;
        RECT 89.265 135.190 91.025 135.420 ;
        RECT 91.355 135.190 93.115 135.420 ;
        RECT 84.805 134.925 85.035 134.985 ;
        RECT 84.740 129.925 85.100 134.925 ;
        RECT 84.805 127.985 85.035 129.925 ;
        RECT 85.425 127.780 86.430 135.190 ;
        RECT 86.895 133.045 87.125 134.985 ;
        RECT 86.830 128.045 87.190 133.045 ;
        RECT 86.895 127.985 87.125 128.045 ;
        RECT 87.520 127.780 88.525 135.190 ;
        RECT 88.985 134.925 89.215 134.985 ;
        RECT 88.920 129.925 89.280 134.925 ;
        RECT 88.985 127.985 89.215 129.925 ;
        RECT 89.635 127.780 90.640 135.190 ;
        RECT 91.075 133.045 91.305 134.985 ;
        RECT 91.010 128.045 91.370 133.045 ;
        RECT 91.075 127.985 91.305 128.045 ;
        RECT 91.665 127.780 92.670 135.190 ;
        RECT 93.165 134.925 93.395 134.985 ;
        RECT 93.100 129.925 93.460 134.925 ;
        RECT 93.165 127.985 93.395 129.925 ;
        RECT 94.205 128.455 95.740 136.005 ;
        RECT 94.225 128.395 95.720 128.455 ;
        RECT 103.760 127.980 104.445 138.930 ;
        RECT 126.985 138.905 128.340 138.930 ;
        RECT 105.270 137.915 110.510 138.145 ;
        RECT 110.840 137.915 121.090 138.145 ;
        RECT 121.420 137.915 126.660 138.145 ;
        RECT 105.270 136.270 105.500 137.915 ;
        RECT 105.175 135.270 105.595 136.270 ;
        RECT 105.270 135.005 105.500 135.270 ;
        RECT 106.275 135.020 109.540 137.915 ;
        RECT 110.560 137.650 110.790 137.710 ;
        RECT 110.495 136.150 110.855 137.650 ;
        RECT 110.560 135.210 110.790 136.150 ;
        RECT 111.705 135.020 114.970 137.915 ;
        RECT 115.850 137.650 116.080 137.915 ;
        RECT 115.755 136.650 116.175 137.650 ;
        RECT 115.850 135.020 116.080 136.650 ;
        RECT 117.055 135.025 120.320 137.915 ;
        RECT 121.140 137.650 121.370 137.710 ;
        RECT 121.075 136.150 121.435 137.650 ;
        RECT 121.140 135.210 121.370 136.150 ;
        RECT 106.275 135.005 110.500 135.020 ;
        RECT 111.705 135.005 116.155 135.020 ;
        RECT 117.055 135.005 121.080 135.025 ;
        RECT 122.220 135.020 125.485 137.915 ;
        RECT 126.430 136.270 126.660 137.915 ;
        RECT 126.335 135.270 126.755 136.270 ;
        RECT 126.430 135.210 126.660 135.270 ;
        RECT 122.220 135.005 126.370 135.020 ;
        RECT 105.270 134.775 110.510 135.005 ;
        RECT 110.840 134.775 121.090 135.005 ;
        RECT 121.420 134.775 126.380 135.005 ;
        RECT 127.680 134.895 128.265 138.905 ;
        RECT 127.700 134.835 128.245 134.895 ;
        RECT 107.200 134.760 110.500 134.775 ;
        RECT 112.490 134.760 116.155 134.775 ;
        RECT 117.780 134.765 121.080 134.775 ;
        RECT 123.070 134.760 126.370 134.775 ;
        RECT 105.515 133.780 129.395 134.280 ;
        RECT 105.530 132.870 127.620 133.370 ;
        RECT 105.270 132.350 105.500 132.355 ;
        RECT 105.270 132.335 108.860 132.350 ;
        RECT 110.850 132.335 114.150 132.350 ;
        RECT 116.140 132.335 119.440 132.350 ;
        RECT 121.430 132.335 124.730 132.350 ;
        RECT 105.270 132.105 110.510 132.335 ;
        RECT 110.840 132.105 121.090 132.335 ;
        RECT 121.420 132.105 126.660 132.335 ;
        RECT 105.270 132.090 109.725 132.105 ;
        RECT 110.850 132.090 114.885 132.105 ;
        RECT 105.270 132.085 105.660 132.090 ;
        RECT 105.270 131.840 105.500 132.085 ;
        RECT 105.175 130.840 105.595 131.840 ;
        RECT 105.270 129.195 105.500 130.840 ;
        RECT 106.460 129.195 109.725 132.090 ;
        RECT 110.560 130.960 110.790 131.900 ;
        RECT 110.495 129.460 110.855 130.960 ;
        RECT 110.560 129.400 110.790 129.460 ;
        RECT 111.620 129.195 114.885 132.090 ;
        RECT 115.850 132.090 120.440 132.105 ;
        RECT 121.430 132.090 125.630 132.105 ;
        RECT 115.850 130.460 116.080 132.090 ;
        RECT 115.755 129.460 116.175 130.460 ;
        RECT 115.850 129.195 116.080 129.460 ;
        RECT 117.175 129.195 120.440 132.090 ;
        RECT 121.140 130.960 121.370 131.900 ;
        RECT 121.075 129.460 121.435 130.960 ;
        RECT 121.140 129.400 121.370 129.460 ;
        RECT 122.365 129.195 125.630 132.090 ;
        RECT 126.430 131.840 126.660 132.105 ;
        RECT 126.335 130.840 126.755 131.840 ;
        RECT 126.430 129.195 126.660 130.840 ;
        RECT 105.270 128.965 110.510 129.195 ;
        RECT 110.840 128.965 121.090 129.195 ;
        RECT 121.420 128.965 126.660 129.195 ;
        RECT 94.140 127.780 94.860 127.825 ;
        RECT 85.085 127.550 94.860 127.780 ;
        RECT 94.140 127.530 94.860 127.550 ;
        RECT 103.760 127.500 126.615 127.980 ;
        RECT 103.780 127.440 126.615 127.500 ;
        RECT 103.925 127.435 126.615 127.440 ;
        RECT 59.030 126.155 71.965 126.900 ;
        RECT 59.050 126.120 71.965 126.155 ;
        RECT 16.565 125.615 51.355 126.120 ;
        RECT 59.050 126.095 59.855 126.120 ;
        RECT 82.970 126.045 93.800 127.285 ;
        RECT 110.570 126.830 110.920 126.860 ;
        RECT 120.935 126.830 121.375 126.860 ;
        RECT 110.570 126.800 121.375 126.830 ;
        RECT 110.550 126.255 121.375 126.800 ;
        RECT 82.970 126.025 84.195 126.045 ;
        RECT 98.460 124.645 99.100 124.740 ;
        RECT 59.330 124.460 60.125 124.520 ;
        RECT 59.310 124.450 60.145 124.460 ;
        RECT 59.310 124.445 60.800 124.450 ;
        RECT 98.410 124.445 99.245 124.645 ;
        RECT 59.310 123.870 99.245 124.445 ;
        RECT 59.310 117.980 60.145 123.870 ;
        RECT 98.410 123.730 99.245 123.870 ;
        RECT 110.550 123.595 110.940 126.255 ;
        RECT 111.475 125.635 113.435 125.865 ;
        RECT 113.765 125.635 115.725 125.865 ;
        RECT 116.055 125.635 118.015 125.865 ;
        RECT 118.345 125.635 120.305 125.865 ;
        RECT 110.570 123.535 110.920 123.595 ;
        RECT 111.195 123.270 111.425 125.475 ;
        RECT 60.990 122.785 70.350 123.015 ;
        RECT 70.680 122.785 89.730 123.015 ;
        RECT 90.060 122.785 99.420 123.015 ;
        RECT 60.710 122.565 60.940 122.625 ;
        RECT 60.615 122.065 61.035 122.565 ;
        RECT 60.710 121.125 60.940 122.065 ;
        RECT 62.090 120.965 69.185 122.785 ;
        RECT 70.400 122.565 70.630 122.625 ;
        RECT 70.335 122.065 70.695 122.565 ;
        RECT 70.400 121.125 70.630 122.065 ;
        RECT 72.260 120.965 79.355 122.785 ;
        RECT 80.090 121.685 80.320 122.785 ;
        RECT 79.995 121.185 80.415 121.685 ;
        RECT 80.090 121.125 80.320 121.185 ;
        RECT 81.405 120.965 88.500 122.785 ;
        RECT 89.780 122.565 90.010 122.625 ;
        RECT 89.715 122.065 90.075 122.565 ;
        RECT 89.780 121.125 90.010 122.065 ;
        RECT 91.255 120.965 98.350 122.785 ;
        RECT 99.470 122.565 99.700 122.625 ;
        RECT 111.015 122.585 111.585 123.270 ;
        RECT 99.375 122.065 99.795 122.565 ;
        RECT 111.195 122.475 111.425 122.585 ;
        RECT 111.855 122.330 112.960 125.635 ;
        RECT 113.485 125.415 113.715 125.475 ;
        RECT 113.420 124.615 113.780 125.415 ;
        RECT 113.485 122.475 113.715 124.615 ;
        RECT 114.150 122.330 115.255 125.635 ;
        RECT 115.775 124.560 116.005 125.475 ;
        RECT 115.610 123.875 116.180 124.560 ;
        RECT 115.775 122.475 116.005 123.875 ;
        RECT 116.465 122.330 117.570 125.635 ;
        RECT 118.065 125.415 118.295 125.475 ;
        RECT 118.000 124.615 118.360 125.415 ;
        RECT 118.065 122.475 118.295 124.615 ;
        RECT 118.735 122.330 119.840 125.635 ;
        RECT 120.355 123.270 120.585 125.475 ;
        RECT 120.190 122.585 120.760 123.270 ;
        RECT 120.355 122.475 120.585 122.585 ;
        RECT 111.855 122.315 113.425 122.330 ;
        RECT 114.150 122.315 115.715 122.330 ;
        RECT 116.465 122.315 118.005 122.330 ;
        RECT 118.735 122.315 120.295 122.330 ;
        RECT 111.475 122.085 113.435 122.315 ;
        RECT 113.765 122.085 115.725 122.315 ;
        RECT 116.055 122.085 118.015 122.315 ;
        RECT 118.345 122.085 120.305 122.315 ;
        RECT 112.325 122.070 113.425 122.085 ;
        RECT 114.615 122.070 115.715 122.085 ;
        RECT 116.905 122.070 118.005 122.085 ;
        RECT 119.195 122.070 120.295 122.085 ;
        RECT 99.470 121.125 99.700 122.065 ;
        RECT 103.630 121.210 120.470 121.710 ;
        RECT 60.990 120.735 99.420 120.965 ;
        RECT 60.710 119.635 60.940 120.575 ;
        RECT 60.615 119.135 61.035 119.635 ;
        RECT 60.710 118.915 60.940 119.135 ;
        RECT 62.110 118.915 69.205 120.735 ;
        RECT 70.400 119.635 70.630 120.575 ;
        RECT 70.335 119.135 70.695 119.635 ;
        RECT 70.400 119.075 70.630 119.135 ;
        RECT 72.240 118.915 79.335 120.735 ;
        RECT 80.090 120.515 80.320 120.575 ;
        RECT 79.995 120.015 80.415 120.515 ;
        RECT 80.090 119.075 80.320 120.015 ;
        RECT 81.405 118.915 88.500 120.735 ;
        RECT 89.780 119.635 90.010 120.575 ;
        RECT 89.715 119.135 90.075 119.635 ;
        RECT 89.780 119.075 90.010 119.135 ;
        RECT 91.255 118.915 98.350 120.735 ;
        RECT 99.470 119.635 99.700 120.575 ;
        RECT 103.580 120.280 120.470 120.780 ;
        RECT 111.485 119.830 112.585 119.845 ;
        RECT 113.775 119.830 114.875 119.845 ;
        RECT 116.065 119.830 117.165 119.845 ;
        RECT 118.355 119.830 119.455 119.845 ;
        RECT 99.375 119.135 99.795 119.635 ;
        RECT 111.475 119.600 113.435 119.830 ;
        RECT 113.765 119.600 115.725 119.830 ;
        RECT 116.055 119.600 118.015 119.830 ;
        RECT 118.345 119.600 120.305 119.830 ;
        RECT 111.485 119.585 112.970 119.600 ;
        RECT 113.775 119.585 115.285 119.600 ;
        RECT 116.065 119.585 117.510 119.600 ;
        RECT 118.355 119.585 119.860 119.600 ;
        RECT 111.195 119.325 111.425 119.440 ;
        RECT 99.470 118.915 99.700 119.135 ;
        RECT 60.710 118.685 70.350 118.915 ;
        RECT 70.680 118.685 80.040 118.915 ;
        RECT 80.370 118.685 89.730 118.915 ;
        RECT 90.060 118.685 99.700 118.915 ;
        RECT 111.020 118.640 111.590 119.325 ;
        RECT 110.525 118.415 110.955 118.475 ;
        RECT 59.300 117.975 60.625 117.980 ;
        RECT 59.300 116.930 99.015 117.975 ;
        RECT 110.505 115.320 110.975 118.415 ;
        RECT 111.195 116.440 111.425 118.640 ;
        RECT 111.865 116.280 112.970 119.585 ;
        RECT 113.485 117.300 113.715 119.440 ;
        RECT 113.420 116.500 113.780 117.300 ;
        RECT 113.485 116.440 113.715 116.500 ;
        RECT 114.180 116.280 115.285 119.585 ;
        RECT 115.775 118.270 116.005 119.440 ;
        RECT 115.605 117.585 116.175 118.270 ;
        RECT 115.775 116.440 116.005 117.585 ;
        RECT 116.405 116.280 117.510 119.585 ;
        RECT 118.065 117.300 118.295 119.440 ;
        RECT 118.000 116.500 118.360 117.300 ;
        RECT 118.065 116.440 118.295 116.500 ;
        RECT 118.755 116.280 119.860 119.585 ;
        RECT 120.355 119.325 120.585 119.440 ;
        RECT 120.180 118.640 120.750 119.325 ;
        RECT 120.355 116.440 120.585 118.640 ;
        RECT 111.475 116.050 113.435 116.280 ;
        RECT 113.765 116.050 115.725 116.280 ;
        RECT 116.055 116.050 118.015 116.280 ;
        RECT 118.345 116.050 120.305 116.280 ;
        RECT 110.300 115.290 111.495 115.320 ;
        RECT 120.935 115.290 121.375 126.255 ;
        RECT 125.985 121.670 126.605 127.435 ;
        RECT 127.120 125.090 127.620 132.870 ;
        RECT 128.895 125.090 129.395 133.780 ;
        RECT 126.935 124.825 127.165 124.885 ;
        RECT 126.870 123.825 127.230 124.825 ;
        RECT 126.935 122.285 127.165 123.825 ;
        RECT 127.575 123.345 127.805 124.885 ;
        RECT 128.715 124.825 128.945 124.885 ;
        RECT 128.650 123.825 129.010 124.825 ;
        RECT 127.510 122.345 127.870 123.345 ;
        RECT 127.575 122.285 127.805 122.345 ;
        RECT 128.715 122.285 128.945 123.825 ;
        RECT 129.355 123.345 129.585 124.885 ;
        RECT 129.290 122.345 129.650 123.345 ;
        RECT 129.355 122.285 129.585 122.345 ;
        RECT 127.205 121.795 127.530 122.085 ;
        RECT 128.995 121.725 129.305 122.080 ;
        RECT 126.005 121.610 126.585 121.670 ;
        RECT 127.510 120.250 127.870 120.415 ;
        RECT 127.325 120.020 129.395 120.250 ;
        RECT 127.605 119.860 127.775 120.020 ;
        RECT 127.135 119.275 127.365 119.860 ;
        RECT 127.070 118.920 127.430 119.275 ;
        RECT 127.135 118.860 127.365 118.920 ;
        RECT 127.575 118.860 127.805 119.860 ;
        RECT 128.915 119.275 129.145 119.860 ;
        RECT 129.355 119.800 129.585 119.860 ;
        RECT 129.290 119.445 129.650 119.800 ;
        RECT 128.850 118.920 129.210 119.275 ;
        RECT 128.915 118.860 129.145 118.920 ;
        RECT 129.355 118.860 129.585 119.445 ;
        RECT 127.325 118.470 129.395 118.700 ;
        RECT 122.995 116.110 130.005 117.530 ;
        RECT 123.025 115.320 123.685 116.110 ;
        RECT 122.680 115.290 123.685 115.320 ;
        RECT 110.300 115.260 123.685 115.290 ;
        RECT 110.280 114.380 123.685 115.260 ;
        RECT 124.485 115.030 125.595 115.040 ;
        RECT 128.655 115.030 129.765 115.035 ;
        RECT 124.475 114.780 126.580 115.030 ;
        RECT 127.670 114.780 129.775 115.030 ;
        RECT 128.655 114.775 129.765 114.780 ;
        RECT 110.280 114.375 117.095 114.380 ;
        RECT 60.235 75.550 61.165 108.560 ;
        RECT 62.390 107.880 63.390 107.975 ;
        RECT 72.675 107.880 73.675 107.945 ;
        RECT 62.330 107.650 66.330 107.880 ;
        RECT 61.940 107.345 62.170 107.600 ;
        RECT 62.390 107.555 63.390 107.650 ;
        RECT 66.490 107.590 66.720 107.600 ;
        RECT 66.475 107.345 66.735 107.590 ;
        RECT 61.940 106.990 66.735 107.345 ;
        RECT 61.940 106.905 66.720 106.990 ;
        RECT 61.940 106.130 62.170 106.905 ;
        RECT 65.270 106.590 66.270 106.665 ;
        RECT 62.330 106.360 66.330 106.590 ;
        RECT 65.270 106.285 66.270 106.360 ;
        RECT 66.490 106.130 66.720 106.905 ;
        RECT 61.940 105.690 66.720 106.130 ;
        RECT 61.940 105.350 62.170 105.690 ;
        RECT 64.150 105.300 64.650 105.365 ;
        RECT 66.490 105.350 66.720 105.690 ;
        RECT 62.330 105.070 66.330 105.300 ;
        RECT 61.940 104.760 62.170 105.020 ;
        RECT 64.150 105.005 64.650 105.070 ;
        RECT 66.490 105.010 66.720 105.020 ;
        RECT 66.475 104.760 66.735 105.010 ;
        RECT 61.940 104.410 66.735 104.760 ;
        RECT 61.940 104.320 66.720 104.410 ;
        RECT 61.940 103.475 62.170 104.320 ;
        RECT 62.390 104.010 63.390 104.075 ;
        RECT 62.330 103.780 66.330 104.010 ;
        RECT 62.390 103.715 63.390 103.780 ;
        RECT 66.490 103.475 66.720 104.320 ;
        RECT 61.940 103.035 66.720 103.475 ;
        RECT 61.940 102.770 62.170 103.035 ;
        RECT 64.150 102.720 64.650 102.785 ;
        RECT 66.490 102.770 66.720 103.035 ;
        RECT 62.330 102.490 66.330 102.720 ;
        RECT 61.940 102.145 62.170 102.440 ;
        RECT 64.150 102.425 64.650 102.490 ;
        RECT 66.490 102.430 66.720 102.440 ;
        RECT 66.475 102.145 66.735 102.430 ;
        RECT 61.940 101.725 66.735 102.145 ;
        RECT 61.940 101.705 66.720 101.725 ;
        RECT 61.940 100.890 62.170 101.705 ;
        RECT 65.270 101.430 66.270 101.505 ;
        RECT 62.330 101.200 66.330 101.430 ;
        RECT 65.270 101.125 66.270 101.200 ;
        RECT 66.490 100.890 66.720 101.705 ;
        RECT 61.940 100.450 66.720 100.890 ;
        RECT 61.940 99.565 62.170 100.450 ;
        RECT 62.390 100.140 63.390 100.235 ;
        RECT 62.330 99.910 66.330 100.140 ;
        RECT 62.390 99.815 63.390 99.910 ;
        RECT 66.490 99.565 66.720 100.450 ;
        RECT 61.940 99.125 66.720 99.565 ;
        RECT 61.940 98.345 62.170 99.125 ;
        RECT 65.270 98.850 66.270 98.925 ;
        RECT 62.330 98.620 66.330 98.850 ;
        RECT 65.270 98.545 66.270 98.620 ;
        RECT 66.490 98.345 66.720 99.125 ;
        RECT 61.940 97.905 66.720 98.345 ;
        RECT 61.940 97.610 62.170 97.905 ;
        RECT 64.150 97.560 64.650 97.625 ;
        RECT 66.490 97.610 66.720 97.905 ;
        RECT 62.330 97.330 66.330 97.560 ;
        RECT 61.940 97.010 62.170 97.280 ;
        RECT 64.150 97.265 64.650 97.330 ;
        RECT 66.490 97.270 66.720 97.280 ;
        RECT 66.475 97.010 66.735 97.270 ;
        RECT 61.940 96.670 66.735 97.010 ;
        RECT 61.940 96.570 66.720 96.670 ;
        RECT 61.940 95.725 62.170 96.570 ;
        RECT 62.390 96.270 63.390 96.330 ;
        RECT 62.330 96.040 66.330 96.270 ;
        RECT 62.390 95.970 63.390 96.040 ;
        RECT 66.490 95.725 66.720 96.570 ;
        RECT 61.940 95.285 66.720 95.725 ;
        RECT 61.940 95.030 62.170 95.285 ;
        RECT 64.150 94.980 64.650 95.045 ;
        RECT 66.490 95.030 66.720 95.285 ;
        RECT 62.330 94.750 66.330 94.980 ;
        RECT 61.940 94.465 62.170 94.700 ;
        RECT 64.150 94.685 64.650 94.750 ;
        RECT 66.490 94.690 66.720 94.700 ;
        RECT 66.475 94.465 66.735 94.690 ;
        RECT 61.940 94.025 66.735 94.465 ;
        RECT 61.940 93.170 62.170 94.025 ;
        RECT 66.475 93.940 66.735 94.025 ;
        RECT 65.270 93.690 66.270 93.765 ;
        RECT 62.330 93.460 66.330 93.690 ;
        RECT 65.270 93.385 66.270 93.460 ;
        RECT 66.490 93.170 66.720 93.940 ;
        RECT 61.940 92.730 66.720 93.170 ;
        RECT 61.940 91.885 62.170 92.730 ;
        RECT 62.390 92.400 63.390 92.495 ;
        RECT 62.330 92.170 66.330 92.400 ;
        RECT 62.390 92.075 63.390 92.170 ;
        RECT 66.490 91.885 66.720 92.730 ;
        RECT 61.940 91.445 66.720 91.885 ;
        RECT 61.940 90.605 62.170 91.445 ;
        RECT 65.270 91.110 66.270 91.185 ;
        RECT 62.330 90.880 66.330 91.110 ;
        RECT 65.270 90.805 66.270 90.880 ;
        RECT 66.490 90.605 66.720 91.445 ;
        RECT 61.940 90.165 66.720 90.605 ;
        RECT 61.940 89.870 62.170 90.165 ;
        RECT 64.150 89.820 64.650 89.885 ;
        RECT 66.490 89.870 66.720 90.165 ;
        RECT 62.330 89.590 66.330 89.820 ;
        RECT 61.940 89.280 62.170 89.540 ;
        RECT 64.150 89.525 64.650 89.590 ;
        RECT 66.490 89.530 66.720 89.540 ;
        RECT 66.475 89.280 66.735 89.530 ;
        RECT 61.940 88.930 66.735 89.280 ;
        RECT 61.940 88.840 66.720 88.930 ;
        RECT 61.940 87.995 62.170 88.840 ;
        RECT 62.390 88.530 63.390 88.595 ;
        RECT 62.330 88.300 66.330 88.530 ;
        RECT 62.390 88.235 63.390 88.300 ;
        RECT 66.490 87.995 66.720 88.840 ;
        RECT 61.940 87.530 66.720 87.995 ;
        RECT 61.940 87.290 62.170 87.530 ;
        RECT 64.150 87.240 64.650 87.305 ;
        RECT 66.490 87.290 66.720 87.530 ;
        RECT 62.330 87.010 66.330 87.240 ;
        RECT 61.940 86.705 62.170 86.960 ;
        RECT 64.150 86.945 64.650 87.010 ;
        RECT 66.490 86.950 66.720 86.960 ;
        RECT 66.475 86.705 66.735 86.950 ;
        RECT 61.940 86.380 66.735 86.705 ;
        RECT 61.940 86.265 66.785 86.380 ;
        RECT 61.940 85.410 62.170 86.265 ;
        RECT 66.425 86.155 66.785 86.265 ;
        RECT 65.270 85.950 66.270 86.025 ;
        RECT 62.330 85.720 66.330 85.950 ;
        RECT 65.270 85.645 66.270 85.720 ;
        RECT 66.490 85.410 66.720 86.155 ;
        RECT 61.940 84.970 66.720 85.410 ;
        RECT 61.940 84.160 62.170 84.970 ;
        RECT 62.390 84.660 63.390 84.755 ;
        RECT 62.330 84.430 66.330 84.660 ;
        RECT 62.390 84.335 63.390 84.430 ;
        RECT 66.490 84.160 66.720 84.970 ;
        RECT 61.940 83.720 66.720 84.160 ;
        RECT 61.940 82.845 62.170 83.720 ;
        RECT 65.270 83.370 66.270 83.445 ;
        RECT 62.330 83.140 66.330 83.370 ;
        RECT 65.270 83.065 66.270 83.140 ;
        RECT 66.490 82.845 66.720 83.720 ;
        RECT 61.940 82.405 66.720 82.845 ;
        RECT 61.940 82.130 62.170 82.405 ;
        RECT 64.150 82.080 64.650 82.145 ;
        RECT 66.490 82.130 66.720 82.405 ;
        RECT 62.330 81.850 66.330 82.080 ;
        RECT 61.940 81.540 62.170 81.800 ;
        RECT 64.150 81.785 64.650 81.850 ;
        RECT 66.490 81.790 66.720 81.800 ;
        RECT 66.475 81.540 66.735 81.790 ;
        RECT 61.940 81.190 66.735 81.540 ;
        RECT 61.940 81.100 66.720 81.190 ;
        RECT 61.940 80.225 62.170 81.100 ;
        RECT 62.390 80.790 63.390 80.855 ;
        RECT 62.330 80.560 66.330 80.790 ;
        RECT 62.390 80.495 63.390 80.560 ;
        RECT 66.490 80.225 66.720 81.100 ;
        RECT 61.940 79.780 66.720 80.225 ;
        RECT 61.940 79.550 62.170 79.780 ;
        RECT 64.150 79.500 64.650 79.565 ;
        RECT 66.490 79.550 66.720 79.780 ;
        RECT 62.330 79.270 66.330 79.500 ;
        RECT 61.940 78.980 62.170 79.220 ;
        RECT 64.150 79.205 64.650 79.270 ;
        RECT 66.490 79.210 66.720 79.220 ;
        RECT 66.475 78.980 66.735 79.210 ;
        RECT 61.940 78.610 66.735 78.980 ;
        RECT 61.940 78.535 66.720 78.610 ;
        RECT 61.940 77.660 62.170 78.535 ;
        RECT 65.270 78.210 66.270 78.285 ;
        RECT 62.330 77.980 66.330 78.210 ;
        RECT 65.270 77.905 66.270 77.980 ;
        RECT 66.490 77.660 66.720 78.535 ;
        RECT 61.940 77.215 66.720 77.660 ;
        RECT 61.940 76.970 62.170 77.215 ;
        RECT 62.390 76.920 63.390 77.015 ;
        RECT 66.490 76.970 66.720 77.215 ;
        RECT 62.330 76.690 66.330 76.920 ;
        RECT 62.390 76.595 63.390 76.690 ;
        RECT 67.605 76.305 67.865 107.830 ;
        RECT 68.330 77.000 68.590 107.830 ;
        RECT 69.735 107.650 73.735 107.880 ;
        RECT 69.345 107.590 69.575 107.600 ;
        RECT 69.330 107.335 69.590 107.590 ;
        RECT 72.675 107.585 73.675 107.650 ;
        RECT 73.895 107.335 74.125 107.600 ;
        RECT 69.330 106.990 74.125 107.335 ;
        RECT 69.345 106.895 74.125 106.990 ;
        RECT 69.345 106.640 69.575 106.895 ;
        RECT 71.300 106.590 71.800 106.655 ;
        RECT 73.895 106.640 74.125 106.895 ;
        RECT 69.735 106.360 73.735 106.590 ;
        RECT 69.345 106.300 69.575 106.310 ;
        RECT 69.330 106.070 69.590 106.300 ;
        RECT 71.300 106.295 71.800 106.360 ;
        RECT 73.895 106.070 74.125 106.310 ;
        RECT 69.330 105.630 74.125 106.070 ;
        RECT 69.330 105.280 69.590 105.630 ;
        RECT 72.675 105.300 73.675 105.375 ;
        RECT 69.345 104.770 69.575 105.280 ;
        RECT 69.735 105.070 73.735 105.300 ;
        RECT 72.675 104.995 73.675 105.070 ;
        RECT 73.895 104.770 74.125 105.630 ;
        RECT 69.345 104.330 74.125 104.770 ;
        RECT 69.345 103.475 69.575 104.330 ;
        RECT 69.795 104.010 70.795 104.105 ;
        RECT 69.735 103.780 73.735 104.010 ;
        RECT 69.795 103.685 70.795 103.780 ;
        RECT 73.895 103.475 74.125 104.330 ;
        RECT 69.345 103.035 74.125 103.475 ;
        RECT 69.345 102.195 69.575 103.035 ;
        RECT 72.675 102.720 73.675 102.795 ;
        RECT 69.735 102.490 73.735 102.720 ;
        RECT 72.675 102.415 73.675 102.490 ;
        RECT 73.895 102.195 74.125 103.035 ;
        RECT 69.345 101.755 74.125 102.195 ;
        RECT 69.345 101.480 69.575 101.755 ;
        RECT 71.300 101.430 71.800 101.495 ;
        RECT 73.895 101.480 74.125 101.755 ;
        RECT 69.735 101.200 73.735 101.430 ;
        RECT 69.345 101.140 69.575 101.150 ;
        RECT 69.330 100.935 69.590 101.140 ;
        RECT 71.300 101.135 71.800 101.200 ;
        RECT 73.895 100.935 74.125 101.150 ;
        RECT 69.330 100.540 74.125 100.935 ;
        RECT 69.345 100.405 74.125 100.540 ;
        RECT 69.345 99.660 69.575 100.405 ;
        RECT 72.675 100.140 73.675 100.205 ;
        RECT 69.735 99.910 73.735 100.140 ;
        RECT 72.675 99.845 73.675 99.910 ;
        RECT 73.895 99.660 74.125 100.405 ;
        RECT 69.345 99.130 74.125 99.660 ;
        RECT 69.345 98.900 69.575 99.130 ;
        RECT 71.300 98.850 71.800 98.915 ;
        RECT 73.895 98.900 74.125 99.130 ;
        RECT 69.735 98.620 73.735 98.850 ;
        RECT 69.345 98.560 69.575 98.570 ;
        RECT 69.330 98.295 69.590 98.560 ;
        RECT 71.300 98.555 71.800 98.620 ;
        RECT 73.895 98.295 74.125 98.570 ;
        RECT 69.330 97.855 74.125 98.295 ;
        RECT 69.330 97.540 69.590 97.855 ;
        RECT 72.675 97.560 73.675 97.635 ;
        RECT 69.345 97.020 69.575 97.540 ;
        RECT 69.735 97.330 73.735 97.560 ;
        RECT 72.675 97.255 73.675 97.330 ;
        RECT 73.895 97.020 74.125 97.855 ;
        RECT 69.345 96.580 74.125 97.020 ;
        RECT 69.345 95.715 69.575 96.580 ;
        RECT 69.795 96.270 70.795 96.365 ;
        RECT 69.735 96.040 73.735 96.270 ;
        RECT 69.795 95.945 70.795 96.040 ;
        RECT 73.895 95.715 74.125 96.580 ;
        RECT 69.345 95.275 74.125 95.715 ;
        RECT 69.345 94.435 69.575 95.275 ;
        RECT 72.675 94.980 73.675 95.055 ;
        RECT 69.735 94.750 73.735 94.980 ;
        RECT 72.675 94.675 73.675 94.750 ;
        RECT 73.895 94.435 74.125 95.275 ;
        RECT 69.345 93.995 74.125 94.435 ;
        RECT 69.345 93.740 69.575 93.995 ;
        RECT 71.295 93.690 71.795 93.755 ;
        RECT 73.895 93.740 74.125 93.995 ;
        RECT 69.735 93.460 73.735 93.690 ;
        RECT 69.345 93.400 69.575 93.410 ;
        RECT 69.330 93.090 69.590 93.400 ;
        RECT 71.295 93.395 71.795 93.460 ;
        RECT 73.895 93.090 74.125 93.410 ;
        RECT 69.330 92.800 74.125 93.090 ;
        RECT 69.345 92.685 74.125 92.800 ;
        RECT 69.345 91.790 69.575 92.685 ;
        RECT 72.675 92.400 73.675 92.465 ;
        RECT 69.735 92.170 73.735 92.400 ;
        RECT 72.675 92.105 73.675 92.170 ;
        RECT 73.895 91.790 74.125 92.685 ;
        RECT 69.345 91.385 74.125 91.790 ;
        RECT 69.345 91.160 69.575 91.385 ;
        RECT 71.300 91.110 71.800 91.175 ;
        RECT 73.895 91.160 74.125 91.385 ;
        RECT 69.735 90.880 73.735 91.110 ;
        RECT 69.345 90.820 69.575 90.830 ;
        RECT 69.330 90.595 69.590 90.820 ;
        RECT 71.300 90.815 71.800 90.880 ;
        RECT 73.895 90.595 74.125 90.830 ;
        RECT 69.330 90.155 74.125 90.595 ;
        RECT 69.330 89.800 69.590 90.155 ;
        RECT 72.675 89.820 73.675 89.895 ;
        RECT 69.345 89.240 69.575 89.800 ;
        RECT 69.735 89.590 73.735 89.820 ;
        RECT 72.675 89.515 73.675 89.590 ;
        RECT 73.895 89.240 74.125 90.155 ;
        RECT 69.345 88.800 74.125 89.240 ;
        RECT 69.345 87.980 69.575 88.800 ;
        RECT 69.795 88.530 70.795 88.625 ;
        RECT 69.735 88.300 73.735 88.530 ;
        RECT 69.795 88.205 70.795 88.300 ;
        RECT 73.895 87.980 74.125 88.800 ;
        RECT 69.345 87.540 74.125 87.980 ;
        RECT 69.345 86.715 69.575 87.540 ;
        RECT 72.675 87.240 73.675 87.315 ;
        RECT 69.735 87.010 73.735 87.240 ;
        RECT 72.675 86.935 73.675 87.010 ;
        RECT 73.895 86.715 74.125 87.540 ;
        RECT 69.345 86.275 74.125 86.715 ;
        RECT 69.345 86.000 69.575 86.275 ;
        RECT 71.300 85.950 71.800 86.015 ;
        RECT 73.895 86.000 74.125 86.275 ;
        RECT 69.735 85.720 73.735 85.950 ;
        RECT 69.345 85.660 69.575 85.670 ;
        RECT 69.330 85.380 69.590 85.660 ;
        RECT 71.300 85.655 71.800 85.720 ;
        RECT 73.895 85.380 74.125 85.670 ;
        RECT 69.330 85.060 74.125 85.380 ;
        RECT 69.345 84.940 74.125 85.060 ;
        RECT 69.345 84.110 69.575 84.940 ;
        RECT 72.675 84.660 73.675 84.725 ;
        RECT 69.735 84.430 73.735 84.660 ;
        RECT 72.675 84.365 73.675 84.430 ;
        RECT 73.895 84.110 74.125 84.940 ;
        RECT 69.345 83.670 74.125 84.110 ;
        RECT 69.345 83.420 69.575 83.670 ;
        RECT 71.300 83.370 71.800 83.435 ;
        RECT 73.895 83.420 74.125 83.670 ;
        RECT 69.735 83.140 73.735 83.370 ;
        RECT 69.345 83.080 69.575 83.090 ;
        RECT 69.330 82.795 69.590 83.080 ;
        RECT 71.300 83.075 71.800 83.140 ;
        RECT 73.895 82.795 74.125 83.090 ;
        RECT 69.330 82.355 74.125 82.795 ;
        RECT 69.330 81.980 69.590 82.355 ;
        RECT 72.675 82.080 73.675 82.155 ;
        RECT 69.345 81.550 69.575 81.980 ;
        RECT 69.735 81.850 73.735 82.080 ;
        RECT 72.675 81.775 73.675 81.850 ;
        RECT 73.895 81.550 74.125 82.355 ;
        RECT 69.345 81.110 74.125 81.550 ;
        RECT 69.345 80.200 69.575 81.110 ;
        RECT 69.795 80.790 70.795 80.885 ;
        RECT 69.735 80.560 73.735 80.790 ;
        RECT 69.795 80.465 70.795 80.560 ;
        RECT 73.895 80.200 74.125 81.110 ;
        RECT 69.345 79.760 74.125 80.200 ;
        RECT 69.345 78.955 69.575 79.760 ;
        RECT 72.670 79.500 73.670 79.575 ;
        RECT 69.735 79.270 73.735 79.500 ;
        RECT 72.670 79.195 73.670 79.270 ;
        RECT 73.895 78.955 74.125 79.760 ;
        RECT 69.345 78.515 74.125 78.955 ;
        RECT 69.345 78.260 69.575 78.515 ;
        RECT 71.300 78.210 71.800 78.275 ;
        RECT 73.895 78.260 74.125 78.515 ;
        RECT 69.735 77.980 73.735 78.210 ;
        RECT 69.345 77.920 69.575 77.930 ;
        RECT 69.330 77.695 69.590 77.920 ;
        RECT 71.300 77.915 71.800 77.980 ;
        RECT 73.895 77.695 74.125 77.930 ;
        RECT 69.330 77.320 74.125 77.695 ;
        RECT 69.345 77.255 74.125 77.320 ;
        RECT 69.345 76.970 69.575 77.255 ;
        RECT 72.675 76.920 73.675 76.985 ;
        RECT 73.895 76.970 74.125 77.255 ;
        RECT 69.735 76.690 73.735 76.920 ;
        RECT 72.675 76.625 73.675 76.690 ;
        RECT 74.940 76.510 75.560 108.340 ;
        RECT 78.650 85.240 79.665 112.395 ;
        RECT 84.415 112.230 85.030 112.295 ;
        RECT 84.355 112.000 85.355 112.230 ;
        RECT 80.480 111.905 80.780 111.970 ;
        RECT 81.060 111.905 81.360 111.970 ;
        RECT 80.420 111.675 81.420 111.905 ;
        RECT 83.920 111.705 84.150 111.975 ;
        RECT 84.415 111.935 85.030 112.000 ;
        RECT 85.560 111.705 85.790 111.950 ;
        RECT 80.030 111.355 80.260 111.625 ;
        RECT 80.480 111.610 80.780 111.675 ;
        RECT 81.060 111.610 81.360 111.675 ;
        RECT 81.580 111.355 81.810 111.625 ;
        RECT 80.030 111.020 81.810 111.355 ;
        RECT 80.030 110.615 80.260 111.020 ;
        RECT 81.580 110.680 81.810 111.020 ;
        RECT 81.060 110.615 81.810 110.680 ;
        RECT 80.030 110.385 81.810 110.615 ;
        RECT 80.030 110.020 80.260 110.385 ;
        RECT 81.060 110.320 81.810 110.385 ;
        RECT 81.580 110.020 81.810 110.320 ;
        RECT 80.030 109.685 81.810 110.020 ;
        RECT 80.030 108.725 80.260 109.685 ;
        RECT 80.480 109.325 80.780 109.390 ;
        RECT 80.420 109.095 81.420 109.325 ;
        RECT 80.480 109.030 80.780 109.095 ;
        RECT 81.580 108.725 81.810 109.685 ;
        RECT 80.030 108.390 81.810 108.725 ;
        RECT 80.030 108.035 80.260 108.390 ;
        RECT 81.580 108.100 81.810 108.390 ;
        RECT 81.060 108.035 81.810 108.100 ;
        RECT 80.030 107.805 81.810 108.035 ;
        RECT 80.030 107.425 80.260 107.805 ;
        RECT 81.060 107.740 81.810 107.805 ;
        RECT 81.580 107.425 81.810 107.740 ;
        RECT 80.030 107.090 81.810 107.425 ;
        RECT 80.030 106.115 80.260 107.090 ;
        RECT 80.480 106.745 80.780 106.810 ;
        RECT 80.420 106.515 81.420 106.745 ;
        RECT 80.480 106.450 80.780 106.515 ;
        RECT 81.580 106.115 81.810 107.090 ;
        RECT 80.030 105.780 81.810 106.115 ;
        RECT 80.030 105.505 80.260 105.780 ;
        RECT 80.480 105.455 80.780 105.520 ;
        RECT 81.580 105.505 81.810 105.780 ;
        RECT 83.920 110.310 85.790 111.705 ;
        RECT 83.920 108.825 84.150 110.310 ;
        RECT 84.680 109.940 85.295 110.005 ;
        RECT 85.560 109.990 85.790 110.310 ;
        RECT 84.355 109.710 85.355 109.940 ;
        RECT 84.680 109.645 85.295 109.710 ;
        RECT 84.415 109.325 85.030 109.390 ;
        RECT 84.355 109.095 85.355 109.325 ;
        RECT 84.415 109.030 85.030 109.095 ;
        RECT 85.560 108.825 85.790 109.045 ;
        RECT 83.920 107.430 85.790 108.825 ;
        RECT 80.420 105.225 81.420 105.455 ;
        RECT 80.030 104.815 80.260 105.175 ;
        RECT 80.480 105.160 80.780 105.225 ;
        RECT 81.580 104.815 81.810 105.175 ;
        RECT 80.030 104.480 81.810 104.815 ;
        RECT 80.030 104.165 80.260 104.480 ;
        RECT 81.580 104.230 81.810 104.480 ;
        RECT 81.060 104.165 81.810 104.230 ;
        RECT 80.030 103.935 81.810 104.165 ;
        RECT 80.030 103.565 80.260 103.935 ;
        RECT 81.060 103.870 81.810 103.935 ;
        RECT 81.580 103.565 81.810 103.870 ;
        RECT 80.030 103.230 81.810 103.565 ;
        RECT 80.030 102.270 80.260 103.230 ;
        RECT 80.480 102.875 80.780 102.940 ;
        RECT 80.420 102.645 81.420 102.875 ;
        RECT 80.480 102.580 80.780 102.645 ;
        RECT 81.580 102.270 81.810 103.230 ;
        RECT 80.030 101.935 81.810 102.270 ;
        RECT 80.030 101.585 80.260 101.935 ;
        RECT 81.580 101.650 81.810 101.935 ;
        RECT 81.060 101.585 81.810 101.650 ;
        RECT 80.030 101.355 81.810 101.585 ;
        RECT 80.030 100.965 80.260 101.355 ;
        RECT 81.060 101.290 81.810 101.355 ;
        RECT 81.580 100.965 81.810 101.290 ;
        RECT 80.030 100.630 81.810 100.965 ;
        RECT 80.030 99.680 80.260 100.630 ;
        RECT 80.480 100.295 80.780 100.360 ;
        RECT 80.420 100.065 81.420 100.295 ;
        RECT 80.480 100.000 80.780 100.065 ;
        RECT 81.580 99.680 81.810 100.630 ;
        RECT 80.030 99.345 81.810 99.680 ;
        RECT 80.030 99.055 80.260 99.345 ;
        RECT 80.480 99.005 80.780 99.070 ;
        RECT 81.580 99.055 81.810 99.345 ;
        RECT 83.920 102.275 84.150 107.430 ;
        RECT 84.675 107.035 85.295 107.100 ;
        RECT 85.560 107.085 85.790 107.430 ;
        RECT 84.355 106.805 85.355 107.035 ;
        RECT 84.675 106.740 85.295 106.805 ;
        RECT 86.620 106.140 87.375 112.535 ;
        RECT 110.280 109.360 112.070 114.375 ;
        RECT 116.615 113.780 118.760 113.830 ;
        RECT 113.270 113.550 118.770 113.780 ;
        RECT 116.615 113.505 118.760 113.550 ;
        RECT 112.880 113.365 113.110 113.500 ;
        RECT 112.805 113.105 113.185 113.365 ;
        RECT 118.930 113.105 119.160 113.500 ;
        RECT 112.805 112.665 119.160 113.105 ;
        RECT 112.880 112.300 119.160 112.665 ;
        RECT 112.880 111.330 113.110 112.300 ;
        RECT 113.280 111.990 115.880 112.035 ;
        RECT 113.270 111.760 118.770 111.990 ;
        RECT 113.280 111.715 115.880 111.760 ;
        RECT 118.930 111.330 119.160 112.300 ;
        RECT 112.880 110.525 119.160 111.330 ;
        RECT 112.880 110.250 113.110 110.525 ;
        RECT 118.930 110.250 119.160 110.525 ;
        RECT 116.615 110.200 118.760 110.250 ;
        RECT 113.270 109.970 118.770 110.200 ;
        RECT 116.615 109.925 118.760 109.970 ;
        RECT 119.725 109.360 120.880 114.380 ;
        RECT 122.680 114.350 123.685 114.380 ;
        RECT 110.280 108.125 120.880 109.360 ;
        RECT 110.300 108.105 120.880 108.125 ;
        RECT 110.300 108.065 111.495 108.105 ;
        RECT 119.725 108.080 120.880 108.105 ;
        RECT 119.745 108.020 120.860 108.080 ;
        RECT 86.600 105.850 87.395 106.140 ;
        RECT 84.415 102.875 84.980 102.940 ;
        RECT 84.355 102.645 85.355 102.875 ;
        RECT 84.415 102.580 84.980 102.645 ;
        RECT 85.560 102.275 85.790 102.595 ;
        RECT 83.920 100.880 85.790 102.275 ;
        RECT 80.420 98.775 81.420 99.005 ;
        RECT 80.030 98.390 80.260 98.725 ;
        RECT 80.480 98.710 80.780 98.775 ;
        RECT 81.580 98.390 81.810 98.725 ;
        RECT 80.030 98.055 81.810 98.390 ;
        RECT 80.030 97.715 80.260 98.055 ;
        RECT 81.580 97.780 81.810 98.055 ;
        RECT 81.060 97.715 81.810 97.780 ;
        RECT 80.030 97.485 81.810 97.715 ;
        RECT 80.030 97.080 80.260 97.485 ;
        RECT 81.060 97.420 81.810 97.485 ;
        RECT 81.580 97.080 81.810 97.420 ;
        RECT 80.030 96.745 81.810 97.080 ;
        RECT 80.030 95.815 80.260 96.745 ;
        RECT 80.480 96.425 80.780 96.490 ;
        RECT 80.420 96.195 81.420 96.425 ;
        RECT 80.480 96.130 80.780 96.195 ;
        RECT 81.580 95.815 81.810 96.745 ;
        RECT 80.030 95.480 81.810 95.815 ;
        RECT 80.030 95.135 80.260 95.480 ;
        RECT 81.580 95.200 81.810 95.480 ;
        RECT 81.060 95.135 81.810 95.200 ;
        RECT 80.030 94.905 81.810 95.135 ;
        RECT 80.030 94.510 80.260 94.905 ;
        RECT 81.060 94.840 81.810 94.905 ;
        RECT 81.580 94.510 81.810 94.840 ;
        RECT 80.030 94.175 81.810 94.510 ;
        RECT 80.030 93.240 80.260 94.175 ;
        RECT 80.480 93.845 80.780 93.910 ;
        RECT 80.420 93.615 81.420 93.845 ;
        RECT 80.480 93.550 80.780 93.615 ;
        RECT 81.580 93.240 81.810 94.175 ;
        RECT 80.030 92.905 81.810 93.240 ;
        RECT 80.030 92.605 80.260 92.905 ;
        RECT 80.480 92.555 80.780 92.620 ;
        RECT 81.580 92.605 81.810 92.905 ;
        RECT 83.920 95.870 84.150 100.880 ;
        RECT 84.680 100.585 85.295 100.650 ;
        RECT 85.560 100.635 85.790 100.880 ;
        RECT 84.355 100.355 85.355 100.585 ;
        RECT 84.680 100.290 85.295 100.355 ;
        RECT 84.415 96.425 84.980 96.490 ;
        RECT 84.355 96.195 85.355 96.425 ;
        RECT 84.415 96.130 84.980 96.195 ;
        RECT 85.560 95.870 85.790 96.145 ;
        RECT 83.920 94.475 85.790 95.870 ;
        RECT 80.420 92.325 81.420 92.555 ;
        RECT 80.030 91.980 80.260 92.275 ;
        RECT 80.480 92.260 80.780 92.325 ;
        RECT 81.580 91.980 81.810 92.275 ;
        RECT 80.030 91.645 81.810 91.980 ;
        RECT 80.030 91.265 80.260 91.645 ;
        RECT 81.580 91.330 81.810 91.645 ;
        RECT 81.060 91.265 81.810 91.330 ;
        RECT 80.030 91.035 81.810 91.265 ;
        RECT 80.030 90.680 80.260 91.035 ;
        RECT 81.060 90.970 81.810 91.035 ;
        RECT 81.580 90.680 81.810 90.970 ;
        RECT 80.030 90.345 81.810 90.680 ;
        RECT 80.030 89.395 80.260 90.345 ;
        RECT 80.480 89.975 80.780 90.040 ;
        RECT 80.420 89.745 81.420 89.975 ;
        RECT 80.480 89.680 80.780 89.745 ;
        RECT 81.580 89.395 81.810 90.345 ;
        RECT 80.030 89.060 81.810 89.395 ;
        RECT 80.030 88.685 80.260 89.060 ;
        RECT 81.580 88.750 81.810 89.060 ;
        RECT 81.060 88.685 81.810 88.750 ;
        RECT 80.030 88.455 81.810 88.685 ;
        RECT 80.030 88.085 80.260 88.455 ;
        RECT 81.060 88.390 81.810 88.455 ;
        RECT 81.580 88.085 81.810 88.390 ;
        RECT 80.030 87.750 81.810 88.085 ;
        RECT 80.030 86.795 80.260 87.750 ;
        RECT 80.480 87.395 80.780 87.460 ;
        RECT 80.420 87.165 81.420 87.395 ;
        RECT 80.480 87.100 80.780 87.165 ;
        RECT 81.580 86.795 81.810 87.750 ;
        RECT 80.030 86.460 81.810 86.795 ;
        RECT 80.030 86.155 80.260 86.460 ;
        RECT 80.480 86.105 80.780 86.170 ;
        RECT 81.580 86.155 81.810 86.460 ;
        RECT 83.920 89.380 84.150 94.475 ;
        RECT 84.680 94.135 85.295 94.200 ;
        RECT 85.560 94.185 85.790 94.475 ;
        RECT 84.355 93.905 85.355 94.135 ;
        RECT 84.680 93.840 85.295 93.905 ;
        RECT 84.415 89.975 84.980 90.040 ;
        RECT 84.355 89.745 85.355 89.975 ;
        RECT 84.415 89.680 84.980 89.745 ;
        RECT 85.560 89.380 85.790 89.695 ;
        RECT 83.920 87.985 85.790 89.380 ;
        RECT 80.420 85.875 81.420 86.105 ;
        RECT 80.480 85.810 80.780 85.875 ;
        RECT 83.920 84.070 84.150 87.985 ;
        RECT 84.680 87.685 85.295 87.750 ;
        RECT 85.560 87.735 85.790 87.985 ;
        RECT 84.355 87.455 85.355 87.685 ;
        RECT 84.680 87.390 85.295 87.455 ;
        RECT 86.620 87.390 87.375 105.850 ;
        RECT 84.415 84.535 85.115 84.630 ;
        RECT 84.355 84.305 85.355 84.535 ;
        RECT 84.415 84.210 85.115 84.305 ;
        RECT 85.560 84.070 85.790 84.255 ;
        RECT 83.920 83.480 85.790 84.070 ;
        RECT 83.920 82.810 84.150 83.480 ;
        RECT 84.595 83.245 85.295 83.310 ;
        RECT 85.560 83.295 85.790 83.480 ;
        RECT 84.355 83.015 85.355 83.245 ;
        RECT 84.595 82.950 85.295 83.015 ;
        RECT 85.560 82.810 85.790 82.965 ;
        RECT 83.920 82.220 85.790 82.810 ;
        RECT 76.670 81.610 81.885 81.630 ;
        RECT 76.610 81.010 81.945 81.610 ;
        RECT 76.670 80.990 81.885 81.010 ;
        RECT 83.920 80.910 84.150 82.220 ;
        RECT 84.415 81.955 85.115 82.050 ;
        RECT 85.560 82.005 85.790 82.220 ;
        RECT 84.355 81.725 85.355 81.955 ;
        RECT 84.415 81.630 85.115 81.725 ;
        RECT 83.920 80.680 84.855 80.910 ;
        RECT 83.920 80.590 84.150 80.680 ;
        RECT 75.745 76.475 76.285 79.230 ;
        RECT 77.875 77.215 80.925 80.265 ;
        RECT 77.875 76.305 78.135 77.215 ;
        RECT 78.835 76.435 81.230 76.455 ;
        RECT 67.605 76.045 78.135 76.305 ;
        RECT 61.545 75.925 62.305 75.945 ;
        RECT 66.495 75.925 67.235 75.945 ;
        RECT 61.485 75.595 62.365 75.925 ;
        RECT 66.435 75.595 67.295 75.925 ;
        RECT 78.775 75.775 81.290 76.435 ;
        RECT 81.690 76.230 82.490 80.475 ;
        RECT 83.815 80.320 84.150 80.590 ;
        RECT 85.060 80.320 85.290 80.630 ;
        RECT 83.815 78.910 85.290 80.320 ;
        RECT 86.050 80.150 86.785 85.200 ;
        RECT 83.815 78.695 84.150 78.910 ;
        RECT 83.920 78.320 84.150 78.695 ;
        RECT 84.415 78.620 84.795 78.685 ;
        RECT 85.060 78.670 85.290 78.910 ;
        RECT 84.355 78.390 84.855 78.620 ;
        RECT 84.415 78.325 84.795 78.390 ;
        RECT 83.815 78.085 84.150 78.320 ;
        RECT 85.060 78.085 85.290 78.340 ;
        RECT 83.815 76.675 85.290 78.085 ;
        RECT 83.815 76.425 84.150 76.675 ;
        RECT 83.920 76.330 84.150 76.425 ;
        RECT 85.060 76.380 85.290 76.675 ;
        RECT 83.920 76.100 84.855 76.330 ;
        RECT 78.835 75.755 81.230 75.775 ;
        RECT 61.545 75.575 62.305 75.595 ;
        RECT 66.495 75.575 67.235 75.595 ;
        RECT 86.060 75.185 86.780 80.150 ;
        RECT 87.115 75.190 87.915 85.205 ;
        RECT 89.490 55.045 128.600 55.550 ;
        RECT 90.140 53.535 127.375 53.765 ;
        RECT 13.410 19.085 14.340 52.095 ;
        RECT 14.720 52.050 15.480 52.070 ;
        RECT 19.670 52.050 20.410 52.070 ;
        RECT 14.660 51.720 15.540 52.050 ;
        RECT 19.610 51.720 20.470 52.050 ;
        RECT 32.010 51.870 34.405 51.890 ;
        RECT 14.720 51.700 15.480 51.720 ;
        RECT 19.670 51.700 20.410 51.720 ;
        RECT 20.780 51.340 31.310 51.600 ;
        RECT 15.565 50.955 16.565 51.050 ;
        RECT 15.505 50.725 19.505 50.955 ;
        RECT 15.115 50.430 15.345 50.675 ;
        RECT 15.565 50.630 16.565 50.725 ;
        RECT 19.665 50.430 19.895 50.675 ;
        RECT 15.115 49.985 19.895 50.430 ;
        RECT 15.115 49.110 15.345 49.985 ;
        RECT 18.445 49.665 19.445 49.740 ;
        RECT 15.505 49.435 19.505 49.665 ;
        RECT 18.445 49.360 19.445 49.435 ;
        RECT 19.665 49.110 19.895 49.985 ;
        RECT 15.115 49.035 19.895 49.110 ;
        RECT 15.115 48.665 19.910 49.035 ;
        RECT 15.115 48.425 15.345 48.665 ;
        RECT 17.325 48.375 17.825 48.440 ;
        RECT 19.650 48.435 19.910 48.665 ;
        RECT 19.665 48.425 19.895 48.435 ;
        RECT 15.505 48.145 19.505 48.375 ;
        RECT 15.115 47.865 15.345 48.095 ;
        RECT 17.325 48.080 17.825 48.145 ;
        RECT 19.665 47.865 19.895 48.095 ;
        RECT 15.115 47.420 19.895 47.865 ;
        RECT 15.115 46.545 15.345 47.420 ;
        RECT 15.565 47.085 16.565 47.150 ;
        RECT 15.505 46.855 19.505 47.085 ;
        RECT 15.565 46.790 16.565 46.855 ;
        RECT 19.665 46.545 19.895 47.420 ;
        RECT 15.115 46.455 19.895 46.545 ;
        RECT 15.115 46.105 19.910 46.455 ;
        RECT 15.115 45.845 15.345 46.105 ;
        RECT 17.325 45.795 17.825 45.860 ;
        RECT 19.650 45.855 19.910 46.105 ;
        RECT 19.665 45.845 19.895 45.855 ;
        RECT 15.505 45.565 19.505 45.795 ;
        RECT 15.115 45.240 15.345 45.515 ;
        RECT 17.325 45.500 17.825 45.565 ;
        RECT 19.665 45.240 19.895 45.515 ;
        RECT 15.115 44.800 19.895 45.240 ;
        RECT 15.115 43.925 15.345 44.800 ;
        RECT 18.445 44.505 19.445 44.580 ;
        RECT 15.505 44.275 19.505 44.505 ;
        RECT 18.445 44.200 19.445 44.275 ;
        RECT 19.665 43.925 19.895 44.800 ;
        RECT 15.115 43.485 19.895 43.925 ;
        RECT 15.115 42.675 15.345 43.485 ;
        RECT 15.565 43.215 16.565 43.310 ;
        RECT 15.505 42.985 19.505 43.215 ;
        RECT 15.565 42.890 16.565 42.985 ;
        RECT 19.665 42.675 19.895 43.485 ;
        RECT 15.115 42.235 19.895 42.675 ;
        RECT 15.115 41.380 15.345 42.235 ;
        RECT 18.445 41.925 19.445 42.000 ;
        RECT 15.505 41.695 19.505 41.925 ;
        RECT 18.445 41.620 19.445 41.695 ;
        RECT 19.665 41.490 19.895 42.235 ;
        RECT 19.600 41.380 19.960 41.490 ;
        RECT 15.115 41.265 19.960 41.380 ;
        RECT 15.115 40.940 19.910 41.265 ;
        RECT 15.115 40.685 15.345 40.940 ;
        RECT 17.325 40.635 17.825 40.700 ;
        RECT 19.650 40.695 19.910 40.940 ;
        RECT 19.665 40.685 19.895 40.695 ;
        RECT 15.505 40.405 19.505 40.635 ;
        RECT 15.115 40.115 15.345 40.355 ;
        RECT 17.325 40.340 17.825 40.405 ;
        RECT 19.665 40.115 19.895 40.355 ;
        RECT 15.115 39.650 19.895 40.115 ;
        RECT 15.115 38.805 15.345 39.650 ;
        RECT 15.565 39.345 16.565 39.410 ;
        RECT 15.505 39.115 19.505 39.345 ;
        RECT 15.565 39.050 16.565 39.115 ;
        RECT 19.665 38.805 19.895 39.650 ;
        RECT 15.115 38.715 19.895 38.805 ;
        RECT 15.115 38.365 19.910 38.715 ;
        RECT 15.115 38.105 15.345 38.365 ;
        RECT 17.325 38.055 17.825 38.120 ;
        RECT 19.650 38.115 19.910 38.365 ;
        RECT 19.665 38.105 19.895 38.115 ;
        RECT 15.505 37.825 19.505 38.055 ;
        RECT 15.115 37.480 15.345 37.775 ;
        RECT 17.325 37.760 17.825 37.825 ;
        RECT 19.665 37.480 19.895 37.775 ;
        RECT 15.115 37.040 19.895 37.480 ;
        RECT 15.115 36.200 15.345 37.040 ;
        RECT 18.445 36.765 19.445 36.840 ;
        RECT 15.505 36.535 19.505 36.765 ;
        RECT 18.445 36.460 19.445 36.535 ;
        RECT 19.665 36.200 19.895 37.040 ;
        RECT 15.115 35.760 19.895 36.200 ;
        RECT 15.115 34.915 15.345 35.760 ;
        RECT 15.565 35.475 16.565 35.570 ;
        RECT 15.505 35.245 19.505 35.475 ;
        RECT 15.565 35.150 16.565 35.245 ;
        RECT 19.665 34.915 19.895 35.760 ;
        RECT 15.115 34.475 19.895 34.915 ;
        RECT 15.115 33.620 15.345 34.475 ;
        RECT 18.445 34.185 19.445 34.260 ;
        RECT 15.505 33.955 19.505 34.185 ;
        RECT 18.445 33.880 19.445 33.955 ;
        RECT 19.665 33.705 19.895 34.475 ;
        RECT 19.650 33.620 19.910 33.705 ;
        RECT 15.115 33.180 19.910 33.620 ;
        RECT 15.115 32.945 15.345 33.180 ;
        RECT 17.325 32.895 17.825 32.960 ;
        RECT 19.650 32.955 19.910 33.180 ;
        RECT 19.665 32.945 19.895 32.955 ;
        RECT 15.505 32.665 19.505 32.895 ;
        RECT 15.115 32.360 15.345 32.615 ;
        RECT 17.325 32.600 17.825 32.665 ;
        RECT 19.665 32.360 19.895 32.615 ;
        RECT 15.115 31.920 19.895 32.360 ;
        RECT 15.115 31.075 15.345 31.920 ;
        RECT 15.565 31.605 16.565 31.675 ;
        RECT 15.505 31.375 19.505 31.605 ;
        RECT 15.565 31.315 16.565 31.375 ;
        RECT 19.665 31.075 19.895 31.920 ;
        RECT 15.115 30.975 19.895 31.075 ;
        RECT 15.115 30.635 19.910 30.975 ;
        RECT 15.115 30.365 15.345 30.635 ;
        RECT 17.325 30.315 17.825 30.380 ;
        RECT 19.650 30.375 19.910 30.635 ;
        RECT 19.665 30.365 19.895 30.375 ;
        RECT 15.505 30.085 19.505 30.315 ;
        RECT 15.115 29.740 15.345 30.035 ;
        RECT 17.325 30.020 17.825 30.085 ;
        RECT 19.665 29.740 19.895 30.035 ;
        RECT 15.115 29.300 19.895 29.740 ;
        RECT 15.115 28.520 15.345 29.300 ;
        RECT 18.445 29.025 19.445 29.100 ;
        RECT 15.505 28.795 19.505 29.025 ;
        RECT 18.445 28.720 19.445 28.795 ;
        RECT 19.665 28.520 19.895 29.300 ;
        RECT 15.115 28.080 19.895 28.520 ;
        RECT 15.115 27.195 15.345 28.080 ;
        RECT 15.565 27.735 16.565 27.830 ;
        RECT 15.505 27.505 19.505 27.735 ;
        RECT 15.565 27.410 16.565 27.505 ;
        RECT 19.665 27.195 19.895 28.080 ;
        RECT 15.115 26.755 19.895 27.195 ;
        RECT 15.115 25.940 15.345 26.755 ;
        RECT 18.445 26.445 19.445 26.520 ;
        RECT 15.505 26.215 19.505 26.445 ;
        RECT 18.445 26.140 19.445 26.215 ;
        RECT 19.665 25.940 19.895 26.755 ;
        RECT 15.115 25.920 19.895 25.940 ;
        RECT 15.115 25.500 19.910 25.920 ;
        RECT 15.115 25.205 15.345 25.500 ;
        RECT 17.325 25.155 17.825 25.220 ;
        RECT 19.650 25.215 19.910 25.500 ;
        RECT 19.665 25.205 19.895 25.215 ;
        RECT 15.505 24.925 19.505 25.155 ;
        RECT 15.115 24.610 15.345 24.875 ;
        RECT 17.325 24.860 17.825 24.925 ;
        RECT 19.665 24.610 19.895 24.875 ;
        RECT 15.115 24.170 19.895 24.610 ;
        RECT 15.115 23.325 15.345 24.170 ;
        RECT 15.565 23.865 16.565 23.930 ;
        RECT 15.505 23.635 19.505 23.865 ;
        RECT 15.565 23.570 16.565 23.635 ;
        RECT 19.665 23.325 19.895 24.170 ;
        RECT 15.115 23.235 19.895 23.325 ;
        RECT 15.115 22.885 19.910 23.235 ;
        RECT 15.115 22.625 15.345 22.885 ;
        RECT 17.325 22.575 17.825 22.640 ;
        RECT 19.650 22.635 19.910 22.885 ;
        RECT 19.665 22.625 19.895 22.635 ;
        RECT 15.505 22.345 19.505 22.575 ;
        RECT 15.115 21.955 15.345 22.295 ;
        RECT 17.325 22.280 17.825 22.345 ;
        RECT 19.665 21.955 19.895 22.295 ;
        RECT 15.115 21.515 19.895 21.955 ;
        RECT 15.115 20.740 15.345 21.515 ;
        RECT 18.445 21.285 19.445 21.360 ;
        RECT 15.505 21.055 19.505 21.285 ;
        RECT 18.445 20.980 19.445 21.055 ;
        RECT 19.665 20.740 19.895 21.515 ;
        RECT 15.115 20.655 19.895 20.740 ;
        RECT 15.115 20.300 19.910 20.655 ;
        RECT 15.115 20.045 15.345 20.300 ;
        RECT 15.565 19.995 16.565 20.090 ;
        RECT 19.650 20.055 19.910 20.300 ;
        RECT 19.665 20.045 19.895 20.055 ;
        RECT 15.505 19.765 19.505 19.995 ;
        RECT 20.780 19.815 21.040 51.340 ;
        RECT 25.850 50.955 26.850 51.020 ;
        RECT 22.910 50.725 26.910 50.955 ;
        RECT 21.505 19.815 21.765 50.645 ;
        RECT 22.520 50.390 22.750 50.675 ;
        RECT 25.850 50.660 26.850 50.725 ;
        RECT 27.070 50.390 27.300 50.675 ;
        RECT 22.520 50.325 27.300 50.390 ;
        RECT 22.505 49.950 27.300 50.325 ;
        RECT 22.505 49.725 22.765 49.950 ;
        RECT 22.520 49.715 22.750 49.725 ;
        RECT 24.475 49.665 24.975 49.730 ;
        RECT 27.070 49.715 27.300 49.950 ;
        RECT 22.910 49.435 26.910 49.665 ;
        RECT 22.520 49.130 22.750 49.385 ;
        RECT 24.475 49.370 24.975 49.435 ;
        RECT 27.070 49.130 27.300 49.385 ;
        RECT 22.520 48.690 27.300 49.130 ;
        RECT 22.520 47.885 22.750 48.690 ;
        RECT 25.845 48.375 26.845 48.450 ;
        RECT 22.910 48.145 26.910 48.375 ;
        RECT 25.845 48.070 26.845 48.145 ;
        RECT 27.070 47.885 27.300 48.690 ;
        RECT 22.520 47.445 27.300 47.885 ;
        RECT 22.520 46.535 22.750 47.445 ;
        RECT 22.970 47.085 23.970 47.180 ;
        RECT 22.910 46.855 26.910 47.085 ;
        RECT 22.970 46.760 23.970 46.855 ;
        RECT 27.070 46.535 27.300 47.445 ;
        RECT 22.520 46.095 27.300 46.535 ;
        RECT 22.520 45.665 22.750 46.095 ;
        RECT 25.850 45.795 26.850 45.870 ;
        RECT 22.505 45.290 22.765 45.665 ;
        RECT 22.910 45.565 26.910 45.795 ;
        RECT 25.850 45.490 26.850 45.565 ;
        RECT 27.070 45.290 27.300 46.095 ;
        RECT 22.505 44.850 27.300 45.290 ;
        RECT 22.505 44.565 22.765 44.850 ;
        RECT 22.520 44.555 22.750 44.565 ;
        RECT 24.475 44.505 24.975 44.570 ;
        RECT 27.070 44.555 27.300 44.850 ;
        RECT 22.910 44.275 26.910 44.505 ;
        RECT 22.520 43.975 22.750 44.225 ;
        RECT 24.475 44.210 24.975 44.275 ;
        RECT 27.070 43.975 27.300 44.225 ;
        RECT 22.520 43.535 27.300 43.975 ;
        RECT 22.520 42.705 22.750 43.535 ;
        RECT 25.850 43.215 26.850 43.280 ;
        RECT 22.910 42.985 26.910 43.215 ;
        RECT 25.850 42.920 26.850 42.985 ;
        RECT 27.070 42.705 27.300 43.535 ;
        RECT 22.520 42.585 27.300 42.705 ;
        RECT 22.505 42.265 27.300 42.585 ;
        RECT 22.505 41.985 22.765 42.265 ;
        RECT 22.520 41.975 22.750 41.985 ;
        RECT 24.475 41.925 24.975 41.990 ;
        RECT 27.070 41.975 27.300 42.265 ;
        RECT 22.910 41.695 26.910 41.925 ;
        RECT 22.520 41.370 22.750 41.645 ;
        RECT 24.475 41.630 24.975 41.695 ;
        RECT 27.070 41.370 27.300 41.645 ;
        RECT 22.520 40.930 27.300 41.370 ;
        RECT 22.520 40.105 22.750 40.930 ;
        RECT 25.850 40.635 26.850 40.710 ;
        RECT 22.910 40.405 26.910 40.635 ;
        RECT 25.850 40.330 26.850 40.405 ;
        RECT 27.070 40.105 27.300 40.930 ;
        RECT 22.520 39.665 27.300 40.105 ;
        RECT 22.520 38.845 22.750 39.665 ;
        RECT 22.970 39.345 23.970 39.440 ;
        RECT 22.910 39.115 26.910 39.345 ;
        RECT 22.970 39.020 23.970 39.115 ;
        RECT 27.070 38.845 27.300 39.665 ;
        RECT 22.520 38.405 27.300 38.845 ;
        RECT 22.520 37.845 22.750 38.405 ;
        RECT 25.850 38.055 26.850 38.130 ;
        RECT 22.505 37.490 22.765 37.845 ;
        RECT 22.910 37.825 26.910 38.055 ;
        RECT 25.850 37.750 26.850 37.825 ;
        RECT 27.070 37.490 27.300 38.405 ;
        RECT 22.505 37.050 27.300 37.490 ;
        RECT 22.505 36.825 22.765 37.050 ;
        RECT 22.520 36.815 22.750 36.825 ;
        RECT 24.475 36.765 24.975 36.830 ;
        RECT 27.070 36.815 27.300 37.050 ;
        RECT 22.910 36.535 26.910 36.765 ;
        RECT 22.520 36.260 22.750 36.485 ;
        RECT 24.475 36.470 24.975 36.535 ;
        RECT 27.070 36.260 27.300 36.485 ;
        RECT 22.520 35.855 27.300 36.260 ;
        RECT 22.520 34.960 22.750 35.855 ;
        RECT 25.850 35.475 26.850 35.540 ;
        RECT 22.910 35.245 26.910 35.475 ;
        RECT 25.850 35.180 26.850 35.245 ;
        RECT 27.070 34.960 27.300 35.855 ;
        RECT 22.520 34.845 27.300 34.960 ;
        RECT 22.505 34.555 27.300 34.845 ;
        RECT 22.505 34.245 22.765 34.555 ;
        RECT 22.520 34.235 22.750 34.245 ;
        RECT 24.470 34.185 24.970 34.250 ;
        RECT 27.070 34.235 27.300 34.555 ;
        RECT 22.910 33.955 26.910 34.185 ;
        RECT 22.520 33.650 22.750 33.905 ;
        RECT 24.470 33.890 24.970 33.955 ;
        RECT 27.070 33.650 27.300 33.905 ;
        RECT 22.520 33.210 27.300 33.650 ;
        RECT 22.520 32.370 22.750 33.210 ;
        RECT 25.850 32.895 26.850 32.970 ;
        RECT 22.910 32.665 26.910 32.895 ;
        RECT 25.850 32.590 26.850 32.665 ;
        RECT 27.070 32.370 27.300 33.210 ;
        RECT 22.520 31.930 27.300 32.370 ;
        RECT 22.520 31.065 22.750 31.930 ;
        RECT 22.970 31.605 23.970 31.700 ;
        RECT 22.910 31.375 26.910 31.605 ;
        RECT 22.970 31.280 23.970 31.375 ;
        RECT 27.070 31.065 27.300 31.930 ;
        RECT 22.520 30.625 27.300 31.065 ;
        RECT 22.520 30.105 22.750 30.625 ;
        RECT 25.850 30.315 26.850 30.390 ;
        RECT 22.505 29.790 22.765 30.105 ;
        RECT 22.910 30.085 26.910 30.315 ;
        RECT 25.850 30.010 26.850 30.085 ;
        RECT 27.070 29.790 27.300 30.625 ;
        RECT 22.505 29.350 27.300 29.790 ;
        RECT 22.505 29.085 22.765 29.350 ;
        RECT 22.520 29.075 22.750 29.085 ;
        RECT 24.475 29.025 24.975 29.090 ;
        RECT 27.070 29.075 27.300 29.350 ;
        RECT 22.910 28.795 26.910 29.025 ;
        RECT 22.520 28.515 22.750 28.745 ;
        RECT 24.475 28.730 24.975 28.795 ;
        RECT 27.070 28.515 27.300 28.745 ;
        RECT 22.520 27.985 27.300 28.515 ;
        RECT 22.520 27.240 22.750 27.985 ;
        RECT 25.850 27.735 26.850 27.800 ;
        RECT 22.910 27.505 26.910 27.735 ;
        RECT 25.850 27.440 26.850 27.505 ;
        RECT 27.070 27.240 27.300 27.985 ;
        RECT 22.520 27.105 27.300 27.240 ;
        RECT 22.505 26.710 27.300 27.105 ;
        RECT 22.505 26.505 22.765 26.710 ;
        RECT 22.520 26.495 22.750 26.505 ;
        RECT 24.475 26.445 24.975 26.510 ;
        RECT 27.070 26.495 27.300 26.710 ;
        RECT 22.910 26.215 26.910 26.445 ;
        RECT 22.520 25.890 22.750 26.165 ;
        RECT 24.475 26.150 24.975 26.215 ;
        RECT 27.070 25.890 27.300 26.165 ;
        RECT 22.520 25.450 27.300 25.890 ;
        RECT 22.520 24.610 22.750 25.450 ;
        RECT 25.850 25.155 26.850 25.230 ;
        RECT 22.910 24.925 26.910 25.155 ;
        RECT 25.850 24.850 26.850 24.925 ;
        RECT 27.070 24.610 27.300 25.450 ;
        RECT 22.520 24.170 27.300 24.610 ;
        RECT 22.520 23.315 22.750 24.170 ;
        RECT 22.970 23.865 23.970 23.960 ;
        RECT 22.910 23.635 26.910 23.865 ;
        RECT 22.970 23.540 23.970 23.635 ;
        RECT 27.070 23.315 27.300 24.170 ;
        RECT 22.520 22.875 27.300 23.315 ;
        RECT 22.520 22.365 22.750 22.875 ;
        RECT 25.850 22.575 26.850 22.650 ;
        RECT 22.505 22.015 22.765 22.365 ;
        RECT 22.910 22.345 26.910 22.575 ;
        RECT 25.850 22.270 26.850 22.345 ;
        RECT 27.070 22.015 27.300 22.875 ;
        RECT 22.505 21.575 27.300 22.015 ;
        RECT 22.505 21.345 22.765 21.575 ;
        RECT 22.520 21.335 22.750 21.345 ;
        RECT 24.475 21.285 24.975 21.350 ;
        RECT 27.070 21.335 27.300 21.575 ;
        RECT 22.910 21.055 26.910 21.285 ;
        RECT 22.520 20.750 22.750 21.005 ;
        RECT 24.475 20.990 24.975 21.055 ;
        RECT 27.070 20.750 27.300 21.005 ;
        RECT 22.520 20.655 27.300 20.750 ;
        RECT 22.505 20.310 27.300 20.655 ;
        RECT 22.505 20.055 22.765 20.310 ;
        RECT 22.520 20.045 22.750 20.055 ;
        RECT 25.850 19.995 26.850 20.060 ;
        RECT 27.070 20.045 27.300 20.310 ;
        RECT 22.910 19.765 26.910 19.995 ;
        RECT 15.565 19.670 16.565 19.765 ;
        RECT 25.850 19.700 26.850 19.765 ;
        RECT 28.115 19.305 28.735 51.135 ;
        RECT 28.920 48.415 29.460 51.170 ;
        RECT 31.050 50.430 31.310 51.340 ;
        RECT 31.950 51.210 34.465 51.870 ;
        RECT 32.010 51.190 34.405 51.210 ;
        RECT 31.050 47.380 34.100 50.430 ;
        RECT 34.865 47.170 35.665 51.415 ;
        RECT 37.095 51.315 38.030 51.545 ;
        RECT 37.095 51.220 37.325 51.315 ;
        RECT 36.990 50.970 37.325 51.220 ;
        RECT 38.235 50.970 38.465 51.265 ;
        RECT 36.990 49.560 38.465 50.970 ;
        RECT 36.990 49.325 37.325 49.560 ;
        RECT 37.095 48.950 37.325 49.325 ;
        RECT 37.590 49.255 37.970 49.320 ;
        RECT 38.235 49.305 38.465 49.560 ;
        RECT 37.530 49.025 38.030 49.255 ;
        RECT 37.590 48.960 37.970 49.025 ;
        RECT 36.990 48.735 37.325 48.950 ;
        RECT 38.235 48.735 38.465 48.975 ;
        RECT 36.990 47.325 38.465 48.735 ;
        RECT 39.235 47.495 39.955 52.460 ;
        RECT 36.990 47.055 37.325 47.325 ;
        RECT 37.095 46.965 37.325 47.055 ;
        RECT 38.235 47.015 38.465 47.325 ;
        RECT 37.095 46.735 38.030 46.965 ;
        RECT 29.845 46.635 35.060 46.655 ;
        RECT 29.785 46.035 35.120 46.635 ;
        RECT 29.845 46.015 35.060 46.035 ;
        RECT 37.095 45.425 37.325 46.735 ;
        RECT 37.590 45.920 38.290 46.015 ;
        RECT 37.530 45.690 38.530 45.920 ;
        RECT 37.590 45.595 38.290 45.690 ;
        RECT 38.735 45.425 38.965 45.640 ;
        RECT 37.095 44.835 38.965 45.425 ;
        RECT 37.095 44.165 37.325 44.835 ;
        RECT 37.770 44.630 38.470 44.695 ;
        RECT 38.735 44.680 38.965 44.835 ;
        RECT 37.530 44.400 38.530 44.630 ;
        RECT 37.770 44.335 38.470 44.400 ;
        RECT 38.735 44.165 38.965 44.350 ;
        RECT 37.095 43.575 38.965 44.165 ;
        RECT 31.825 14.755 32.840 41.910 ;
        RECT 33.655 41.275 33.955 41.340 ;
        RECT 33.595 41.045 34.595 41.275 ;
        RECT 33.205 40.690 33.435 40.995 ;
        RECT 33.655 40.980 33.955 41.045 ;
        RECT 34.755 40.690 34.985 40.995 ;
        RECT 33.205 40.355 34.985 40.690 ;
        RECT 33.205 39.400 33.435 40.355 ;
        RECT 33.655 39.985 33.955 40.050 ;
        RECT 33.595 39.755 34.595 39.985 ;
        RECT 33.655 39.690 33.955 39.755 ;
        RECT 34.755 39.400 34.985 40.355 ;
        RECT 33.205 39.065 34.985 39.400 ;
        RECT 33.205 38.695 33.435 39.065 ;
        RECT 34.755 38.760 34.985 39.065 ;
        RECT 34.235 38.695 34.985 38.760 ;
        RECT 33.205 38.465 34.985 38.695 ;
        RECT 33.205 38.090 33.435 38.465 ;
        RECT 34.235 38.400 34.985 38.465 ;
        RECT 34.755 38.090 34.985 38.400 ;
        RECT 33.205 37.755 34.985 38.090 ;
        RECT 33.205 36.805 33.435 37.755 ;
        RECT 33.655 37.405 33.955 37.470 ;
        RECT 33.595 37.175 34.595 37.405 ;
        RECT 33.655 37.110 33.955 37.175 ;
        RECT 34.755 36.805 34.985 37.755 ;
        RECT 33.205 36.470 34.985 36.805 ;
        RECT 33.205 36.115 33.435 36.470 ;
        RECT 34.755 36.180 34.985 36.470 ;
        RECT 34.235 36.115 34.985 36.180 ;
        RECT 33.205 35.885 34.985 36.115 ;
        RECT 33.205 35.505 33.435 35.885 ;
        RECT 34.235 35.820 34.985 35.885 ;
        RECT 34.755 35.505 34.985 35.820 ;
        RECT 33.205 35.170 34.985 35.505 ;
        RECT 33.205 34.875 33.435 35.170 ;
        RECT 33.655 34.825 33.955 34.890 ;
        RECT 34.755 34.875 34.985 35.170 ;
        RECT 37.095 39.165 37.325 43.575 ;
        RECT 37.590 43.340 38.290 43.435 ;
        RECT 38.735 43.390 38.965 43.575 ;
        RECT 37.530 43.110 38.530 43.340 ;
        RECT 37.590 43.015 38.290 43.110 ;
        RECT 39.225 42.445 39.960 47.495 ;
        RECT 40.290 42.440 41.090 52.455 ;
        RECT 90.140 51.525 91.140 53.535 ;
        RECT 90.140 46.370 90.570 51.525 ;
        RECT 92.025 51.325 108.220 53.535 ;
        RECT 109.135 53.270 109.365 53.330 ;
        RECT 109.065 51.590 109.435 53.270 ;
        RECT 109.135 51.530 109.365 51.590 ;
        RECT 110.335 51.325 126.530 53.535 ;
        RECT 127.355 51.535 128.365 53.335 ;
        RECT 127.425 51.530 127.655 51.535 ;
        RECT 91.125 51.095 109.085 51.325 ;
        RECT 109.415 51.095 127.375 51.325 ;
        RECT 90.710 49.085 91.140 50.890 ;
        RECT 92.025 48.885 108.220 51.095 ;
        RECT 109.135 50.830 109.365 50.890 ;
        RECT 109.065 49.150 109.435 50.830 ;
        RECT 109.135 49.090 109.365 49.150 ;
        RECT 110.335 48.885 126.530 51.095 ;
        RECT 127.365 48.885 127.795 50.890 ;
        RECT 91.125 48.655 127.795 48.885 ;
        RECT 127.935 47.295 128.365 51.535 ;
        RECT 90.710 47.290 129.505 47.295 ;
        RECT 132.440 47.290 133.440 47.295 ;
        RECT 90.710 46.795 133.440 47.290 ;
        RECT 129.430 46.790 133.440 46.795 ;
        RECT 132.440 46.490 133.440 46.790 ;
        RECT 90.140 45.870 127.845 46.370 ;
        RECT 97.175 44.130 109.135 44.360 ;
        RECT 109.465 44.130 121.425 44.360 ;
        RECT 96.895 43.910 97.125 43.970 ;
        RECT 37.855 39.695 38.470 39.760 ;
        RECT 37.530 39.465 38.530 39.695 ;
        RECT 37.855 39.400 38.470 39.465 ;
        RECT 38.735 39.165 38.965 39.415 ;
        RECT 37.095 37.770 38.965 39.165 ;
        RECT 33.595 34.595 34.595 34.825 ;
        RECT 33.205 34.245 33.435 34.545 ;
        RECT 33.655 34.530 33.955 34.595 ;
        RECT 34.755 34.245 34.985 34.545 ;
        RECT 33.205 33.910 34.985 34.245 ;
        RECT 33.205 32.975 33.435 33.910 ;
        RECT 33.655 33.535 33.955 33.600 ;
        RECT 33.595 33.305 34.595 33.535 ;
        RECT 33.655 33.240 33.955 33.305 ;
        RECT 34.755 32.975 34.985 33.910 ;
        RECT 33.205 32.640 34.985 32.975 ;
        RECT 33.205 32.245 33.435 32.640 ;
        RECT 34.755 32.310 34.985 32.640 ;
        RECT 34.235 32.245 34.985 32.310 ;
        RECT 33.205 32.015 34.985 32.245 ;
        RECT 33.205 31.670 33.435 32.015 ;
        RECT 34.235 31.950 34.985 32.015 ;
        RECT 34.755 31.670 34.985 31.950 ;
        RECT 33.205 31.335 34.985 31.670 ;
        RECT 33.205 30.405 33.435 31.335 ;
        RECT 33.655 30.955 33.955 31.020 ;
        RECT 33.595 30.725 34.595 30.955 ;
        RECT 33.655 30.660 33.955 30.725 ;
        RECT 34.755 30.405 34.985 31.335 ;
        RECT 33.205 30.070 34.985 30.405 ;
        RECT 33.205 29.665 33.435 30.070 ;
        RECT 34.755 29.730 34.985 30.070 ;
        RECT 34.235 29.665 34.985 29.730 ;
        RECT 33.205 29.435 34.985 29.665 ;
        RECT 33.205 29.095 33.435 29.435 ;
        RECT 34.235 29.370 34.985 29.435 ;
        RECT 34.755 29.095 34.985 29.370 ;
        RECT 33.205 28.760 34.985 29.095 ;
        RECT 33.205 28.425 33.435 28.760 ;
        RECT 33.655 28.375 33.955 28.440 ;
        RECT 34.755 28.425 34.985 28.760 ;
        RECT 37.095 32.675 37.325 37.770 ;
        RECT 37.590 37.405 38.155 37.470 ;
        RECT 38.735 37.455 38.965 37.770 ;
        RECT 37.530 37.175 38.530 37.405 ;
        RECT 37.590 37.110 38.155 37.175 ;
        RECT 37.855 33.245 38.470 33.310 ;
        RECT 37.530 33.015 38.530 33.245 ;
        RECT 37.855 32.950 38.470 33.015 ;
        RECT 38.735 32.675 38.965 32.965 ;
        RECT 37.095 31.280 38.965 32.675 ;
        RECT 33.595 28.145 34.595 28.375 ;
        RECT 33.205 27.805 33.435 28.095 ;
        RECT 33.655 28.080 33.955 28.145 ;
        RECT 34.755 27.805 34.985 28.095 ;
        RECT 33.205 27.470 34.985 27.805 ;
        RECT 33.205 26.520 33.435 27.470 ;
        RECT 33.655 27.085 33.955 27.150 ;
        RECT 33.595 26.855 34.595 27.085 ;
        RECT 33.655 26.790 33.955 26.855 ;
        RECT 34.755 26.520 34.985 27.470 ;
        RECT 33.205 26.185 34.985 26.520 ;
        RECT 33.205 25.795 33.435 26.185 ;
        RECT 34.755 25.860 34.985 26.185 ;
        RECT 34.235 25.795 34.985 25.860 ;
        RECT 33.205 25.565 34.985 25.795 ;
        RECT 33.205 25.215 33.435 25.565 ;
        RECT 34.235 25.500 34.985 25.565 ;
        RECT 34.755 25.215 34.985 25.500 ;
        RECT 33.205 24.880 34.985 25.215 ;
        RECT 33.205 23.920 33.435 24.880 ;
        RECT 33.655 24.505 33.955 24.570 ;
        RECT 33.595 24.275 34.595 24.505 ;
        RECT 33.655 24.210 33.955 24.275 ;
        RECT 34.755 23.920 34.985 24.880 ;
        RECT 33.205 23.585 34.985 23.920 ;
        RECT 33.205 23.215 33.435 23.585 ;
        RECT 34.755 23.280 34.985 23.585 ;
        RECT 34.235 23.215 34.985 23.280 ;
        RECT 33.205 22.985 34.985 23.215 ;
        RECT 33.205 22.670 33.435 22.985 ;
        RECT 34.235 22.920 34.985 22.985 ;
        RECT 34.755 22.670 34.985 22.920 ;
        RECT 33.205 22.335 34.985 22.670 ;
        RECT 33.205 21.975 33.435 22.335 ;
        RECT 33.655 21.925 33.955 21.990 ;
        RECT 34.755 21.975 34.985 22.335 ;
        RECT 37.095 26.270 37.325 31.280 ;
        RECT 37.590 30.955 38.155 31.020 ;
        RECT 38.735 31.005 38.965 31.280 ;
        RECT 37.530 30.725 38.530 30.955 ;
        RECT 37.590 30.660 38.155 30.725 ;
        RECT 37.855 26.795 38.470 26.860 ;
        RECT 37.530 26.565 38.530 26.795 ;
        RECT 37.855 26.500 38.470 26.565 ;
        RECT 38.735 26.270 38.965 26.515 ;
        RECT 37.095 24.875 38.965 26.270 ;
        RECT 33.595 21.695 34.595 21.925 ;
        RECT 33.205 21.370 33.435 21.645 ;
        RECT 33.655 21.630 33.955 21.695 ;
        RECT 34.755 21.370 34.985 21.645 ;
        RECT 33.205 21.035 34.985 21.370 ;
        RECT 33.205 20.060 33.435 21.035 ;
        RECT 33.655 20.635 33.955 20.700 ;
        RECT 33.595 20.405 34.595 20.635 ;
        RECT 33.655 20.340 33.955 20.405 ;
        RECT 34.755 20.060 34.985 21.035 ;
        RECT 33.205 19.725 34.985 20.060 ;
        RECT 33.205 19.345 33.435 19.725 ;
        RECT 34.755 19.410 34.985 19.725 ;
        RECT 34.235 19.345 34.985 19.410 ;
        RECT 33.205 19.115 34.985 19.345 ;
        RECT 33.205 18.760 33.435 19.115 ;
        RECT 34.235 19.050 34.985 19.115 ;
        RECT 34.755 18.760 34.985 19.050 ;
        RECT 33.205 18.425 34.985 18.760 ;
        RECT 33.205 17.465 33.435 18.425 ;
        RECT 33.655 18.055 33.955 18.120 ;
        RECT 33.595 17.825 34.595 18.055 ;
        RECT 33.655 17.760 33.955 17.825 ;
        RECT 34.755 17.465 34.985 18.425 ;
        RECT 33.205 17.130 34.985 17.465 ;
        RECT 33.205 16.765 33.435 17.130 ;
        RECT 34.755 16.830 34.985 17.130 ;
        RECT 34.235 16.765 34.985 16.830 ;
        RECT 33.205 16.535 34.985 16.765 ;
        RECT 33.205 16.130 33.435 16.535 ;
        RECT 34.235 16.470 34.985 16.535 ;
        RECT 34.755 16.130 34.985 16.470 ;
        RECT 33.205 15.795 34.985 16.130 ;
        RECT 33.205 15.525 33.435 15.795 ;
        RECT 33.655 15.475 33.955 15.540 ;
        RECT 34.235 15.475 34.535 15.540 ;
        RECT 34.755 15.525 34.985 15.795 ;
        RECT 37.095 19.720 37.325 24.875 ;
        RECT 37.590 24.505 38.155 24.570 ;
        RECT 38.735 24.555 38.965 24.875 ;
        RECT 37.530 24.275 38.530 24.505 ;
        RECT 37.590 24.210 38.155 24.275 ;
        RECT 39.795 21.300 40.550 39.760 ;
        RECT 96.655 38.240 97.185 43.910 ;
        RECT 96.895 37.970 97.125 38.240 ;
        RECT 100.415 37.840 105.840 44.130 ;
        RECT 109.185 39.785 109.415 43.970 ;
        RECT 109.125 38.190 109.485 39.785 ;
        RECT 109.185 37.970 109.415 38.190 ;
        RECT 112.935 37.840 118.370 44.130 ;
        RECT 121.475 43.910 121.705 43.970 ;
        RECT 121.415 38.305 121.945 43.910 ;
        RECT 121.475 37.970 121.705 38.305 ;
        RECT 97.205 37.810 109.125 37.840 ;
        RECT 109.475 37.810 121.415 37.840 ;
        RECT 97.175 37.580 109.135 37.810 ;
        RECT 109.465 37.580 121.425 37.810 ;
        RECT 97.205 37.555 109.125 37.580 ;
        RECT 109.475 37.555 121.415 37.580 ;
        RECT 97.255 36.875 110.570 37.270 ;
        RECT 90.240 36.375 93.220 36.430 ;
        RECT 90.230 36.145 93.230 36.375 ;
        RECT 89.840 35.100 90.070 36.095 ;
        RECT 93.390 35.190 93.685 36.095 ;
        RECT 108.020 35.340 121.365 35.785 ;
        RECT 93.330 35.100 93.690 35.190 ;
        RECT 89.840 32.115 93.690 35.100 ;
        RECT 97.180 34.985 109.120 35.015 ;
        RECT 109.470 34.985 121.410 35.010 ;
        RECT 97.170 34.755 109.130 34.985 ;
        RECT 109.460 34.755 121.420 34.985 ;
        RECT 97.180 34.730 109.120 34.755 ;
        RECT 96.890 34.535 97.120 34.595 ;
        RECT 89.840 31.135 90.070 32.115 ;
        RECT 93.330 31.195 93.690 32.115 ;
        RECT 93.390 31.135 93.685 31.195 ;
        RECT 90.230 30.855 93.230 31.085 ;
        RECT 96.125 28.830 97.180 34.535 ;
        RECT 96.890 28.595 97.120 28.830 ;
        RECT 100.390 28.440 105.825 34.730 ;
        RECT 109.470 34.725 121.410 34.755 ;
        RECT 109.180 34.380 109.410 34.595 ;
        RECT 109.120 32.785 109.480 34.380 ;
        RECT 109.180 28.595 109.410 32.785 ;
        RECT 89.100 27.835 91.985 28.365 ;
        RECT 97.170 28.180 109.130 28.440 ;
        RECT 109.470 28.435 111.970 28.445 ;
        RECT 112.890 28.435 118.325 34.725 ;
        RECT 121.470 34.535 121.700 34.595 ;
        RECT 121.405 29.175 122.265 34.535 ;
        RECT 121.470 28.595 121.700 29.175 ;
        RECT 109.460 28.205 121.420 28.435 ;
        RECT 109.470 28.185 111.970 28.205 ;
        RECT 89.110 26.685 123.900 27.190 ;
        RECT 39.775 21.010 40.570 21.300 ;
        RECT 37.850 20.345 38.470 20.410 ;
        RECT 37.530 20.115 38.530 20.345 ;
        RECT 37.850 20.050 38.470 20.115 ;
        RECT 38.735 19.720 38.965 20.065 ;
        RECT 37.095 18.325 38.965 19.720 ;
        RECT 37.095 16.840 37.325 18.325 ;
        RECT 37.590 18.055 38.205 18.120 ;
        RECT 38.735 18.105 38.965 18.325 ;
        RECT 37.530 17.825 38.530 18.055 ;
        RECT 37.590 17.760 38.205 17.825 ;
        RECT 37.855 17.440 38.470 17.505 ;
        RECT 37.530 17.210 38.530 17.440 ;
        RECT 37.855 17.145 38.470 17.210 ;
        RECT 38.735 16.840 38.965 17.160 ;
        RECT 33.595 15.245 34.595 15.475 ;
        RECT 37.095 15.445 38.965 16.840 ;
        RECT 33.655 15.180 33.955 15.245 ;
        RECT 34.235 15.180 34.535 15.245 ;
        RECT 37.095 15.175 37.325 15.445 ;
        RECT 37.590 15.150 38.205 15.215 ;
        RECT 38.735 15.200 38.965 15.445 ;
        RECT 37.530 14.920 38.530 15.150 ;
        RECT 37.590 14.855 38.205 14.920 ;
        RECT 39.795 14.615 40.550 21.010 ;
      LAYER met2 ;
        RECT 58.555 163.995 71.960 165.110 ;
        RECT 58.555 163.990 59.825 163.995 ;
        RECT 58.560 155.965 59.825 163.990 ;
        RECT 62.785 162.130 76.190 162.630 ;
        RECT 62.785 159.530 63.145 162.130 ;
        RECT 67.165 159.530 67.525 162.130 ;
        RECT 56.190 155.955 59.825 155.965 ;
        RECT 16.085 153.955 59.825 155.955 ;
        RECT 18.115 146.240 18.545 149.820 ;
        RECT 36.570 148.030 36.840 153.955 ;
        RECT 56.190 153.950 59.825 153.955 ;
        RECT 18.115 145.720 19.710 146.240 ;
        RECT 22.205 145.725 24.010 146.225 ;
        RECT 47.525 145.725 49.350 146.225 ;
        RECT 17.745 135.035 20.625 135.460 ;
        RECT 20.835 134.165 21.095 134.170 ;
        RECT 20.820 130.075 21.110 134.165 ;
        RECT 23.580 133.515 24.010 145.725 ;
        RECT 24.160 144.800 26.090 145.300 ;
        RECT 24.160 139.950 24.590 144.800 ;
        RECT 48.920 139.950 49.350 145.725 ;
        RECT 54.870 145.300 55.300 149.820 ;
        RECT 59.000 146.955 59.825 153.950 ;
        RECT 64.995 153.835 65.315 158.935 ;
        RECT 60.610 147.650 60.930 152.750 ;
        RECT 69.375 147.650 69.695 152.750 ;
        RECT 61.000 147.140 62.400 147.500 ;
        RECT 63.190 147.140 64.590 147.500 ;
        RECT 65.380 147.140 66.780 147.500 ;
        RECT 67.570 147.140 68.970 147.500 ;
        RECT 61.000 145.675 61.500 147.140 ;
        RECT 49.500 144.800 51.370 145.300 ;
        RECT 53.195 144.800 55.300 145.300 ;
        RECT 36.610 137.020 36.890 138.830 ;
        RECT 24.710 135.845 25.760 136.820 ;
        RECT 35.475 133.610 36.525 134.655 ;
        RECT 36.975 133.605 38.025 136.260 ;
        RECT 47.770 134.280 48.820 136.820 ;
        RECT 49.500 133.515 49.930 144.800 ;
        RECT 62.240 143.255 62.740 144.730 ;
        RECT 63.190 144.130 63.690 147.140 ;
        RECT 64.430 143.255 64.930 146.275 ;
        RECT 65.380 144.130 65.880 147.140 ;
        RECT 66.620 143.255 67.120 146.275 ;
        RECT 67.570 145.675 68.070 147.140 ;
        RECT 68.810 143.255 69.310 144.730 ;
        RECT 23.580 130.645 24.585 133.515 ;
        RECT 36.605 131.615 36.895 133.410 ;
        RECT 23.580 127.760 24.595 130.645 ;
        RECT 48.910 128.055 49.930 133.515 ;
        RECT 15.075 127.595 15.565 127.645 ;
        RECT 15.075 126.140 19.985 127.595 ;
        RECT 24.685 127.045 27.085 127.435 ;
        RECT 36.975 127.055 39.375 127.445 ;
        RECT 59.085 127.085 59.825 142.965 ;
        RECT 61.340 142.895 62.740 143.255 ;
        RECT 63.530 142.895 64.930 143.255 ;
        RECT 65.720 142.895 67.120 143.255 ;
        RECT 67.910 142.895 69.310 143.255 ;
        RECT 60.615 137.645 60.935 142.745 ;
        RECT 69.375 137.645 69.695 142.745 ;
        RECT 64.995 131.845 65.315 136.945 ;
        RECT 75.690 134.975 76.190 162.130 ;
        RECT 76.645 145.675 78.105 146.275 ;
        RECT 93.695 140.835 103.755 140.855 ;
        RECT 135.140 140.850 136.630 140.905 ;
        RECT 128.445 140.845 136.630 140.850 ;
        RECT 128.210 140.840 136.630 140.845 ;
        RECT 127.015 140.835 136.630 140.840 ;
        RECT 93.695 138.920 136.630 140.835 ;
        RECT 93.695 138.915 128.310 138.920 ;
        RECT 93.695 138.910 127.520 138.915 ;
        RECT 93.695 138.905 104.535 138.910 ;
        RECT 93.695 137.540 95.690 138.905 ;
        RECT 103.460 138.765 104.535 138.905 ;
        RECT 77.375 135.985 95.690 137.540 ;
        RECT 75.690 134.475 93.410 134.975 ;
        RECT 62.785 130.865 69.785 130.870 ;
        RECT 75.690 130.865 76.190 134.475 ;
        RECT 62.785 130.370 76.190 130.865 ;
        RECT 62.785 127.765 63.145 130.370 ;
        RECT 67.160 127.765 67.520 130.370 ;
        RECT 69.145 130.365 76.190 130.370 ;
        RECT 84.790 129.875 85.050 134.475 ;
        RECT 86.880 127.305 87.140 133.095 ;
        RECT 88.970 129.875 89.230 134.475 ;
        RECT 91.060 127.305 91.320 133.095 ;
        RECT 93.150 129.875 93.410 134.475 ;
        RECT 94.255 128.405 95.690 135.985 ;
        RECT 103.810 128.000 104.395 138.765 ;
        RECT 105.225 135.220 105.545 136.320 ;
        RECT 110.545 136.100 110.805 138.910 ;
        RECT 115.805 136.600 116.125 137.700 ;
        RECT 121.125 136.100 121.385 138.910 ;
        RECT 126.385 135.220 126.705 136.320 ;
        RECT 107.250 134.710 110.450 135.070 ;
        RECT 112.540 134.710 115.740 135.070 ;
        RECT 117.830 134.715 121.030 135.075 ;
        RECT 109.950 133.730 110.450 134.710 ;
        RECT 105.610 132.400 106.110 133.420 ;
        RECT 110.900 132.400 111.400 134.330 ;
        RECT 115.240 132.820 115.740 134.710 ;
        RECT 116.190 132.400 116.690 134.330 ;
        RECT 120.530 132.820 121.030 134.715 ;
        RECT 123.120 134.710 126.320 135.070 ;
        RECT 127.730 134.845 128.215 138.915 ;
        RECT 135.140 138.870 136.630 138.920 ;
        RECT 125.820 133.730 126.320 134.710 ;
        RECT 121.480 132.400 121.980 133.420 ;
        RECT 105.610 132.040 108.810 132.400 ;
        RECT 110.900 132.040 114.100 132.400 ;
        RECT 116.190 132.040 119.390 132.400 ;
        RECT 121.480 132.040 124.680 132.400 ;
        RECT 105.225 130.790 105.545 131.890 ;
        RECT 110.545 128.000 110.805 131.010 ;
        RECT 115.805 129.410 116.125 130.510 ;
        RECT 121.125 128.000 121.385 131.010 ;
        RECT 126.385 130.790 126.705 131.890 ;
        RECT 94.190 127.480 102.250 127.875 ;
        RECT 59.080 126.920 59.825 127.085 ;
        RECT 15.075 125.595 51.295 126.140 ;
        RECT 59.080 126.105 71.905 126.920 ;
        RECT 59.645 126.100 71.905 126.105 ;
        RECT 83.425 126.025 93.740 127.305 ;
        RECT 15.075 125.545 15.565 125.595 ;
        RECT 49.250 124.475 51.295 125.595 ;
        RECT 59.360 124.475 60.095 124.510 ;
        RECT 49.235 124.470 60.095 124.475 ;
        RECT 49.235 124.465 60.740 124.470 ;
        RECT 98.460 124.465 99.195 124.695 ;
        RECT 49.235 123.850 99.195 124.465 ;
        RECT 49.235 122.790 60.095 123.850 ;
        RECT 45.645 118.000 46.915 118.050 ;
        RECT 59.360 118.020 60.095 122.790 ;
        RECT 60.665 122.015 60.985 122.615 ;
        RECT 70.385 122.015 70.645 123.850 ;
        RECT 89.765 122.015 90.025 123.850 ;
        RECT 98.460 123.680 99.195 123.850 ;
        RECT 99.425 122.015 99.745 122.615 ;
        RECT 80.045 121.135 80.365 121.735 ;
        RECT 80.045 119.965 80.365 120.565 ;
        RECT 60.665 119.085 60.985 119.685 ;
        RECT 70.385 118.020 70.645 119.685 ;
        RECT 89.765 118.020 90.025 119.685 ;
        RECT 99.425 119.085 99.745 119.685 ;
        RECT 59.350 118.000 96.625 118.020 ;
        RECT 45.645 117.995 96.625 118.000 ;
        RECT 99.295 117.995 100.215 118.045 ;
        RECT 45.645 116.910 100.260 117.995 ;
        RECT 45.645 116.860 46.915 116.910 ;
        RECT 59.350 116.905 96.625 116.910 ;
        RECT 60.210 107.570 61.185 116.905 ;
        RECT 99.295 116.860 100.215 116.910 ;
        RECT 64.100 108.695 71.850 109.295 ;
        RECT 62.340 107.605 63.440 107.925 ;
        RECT 57.630 106.705 58.415 106.755 ;
        RECT 60.215 106.705 61.185 107.570 ;
        RECT 57.630 104.840 61.185 106.705 ;
        RECT 57.630 104.790 58.415 104.840 ;
        RECT 60.215 104.025 61.185 104.840 ;
        RECT 64.100 104.670 64.700 108.695 ;
        RECT 67.555 107.540 67.915 107.780 ;
        RECT 66.425 107.280 67.915 107.540 ;
        RECT 68.280 107.540 68.640 107.780 ;
        RECT 68.280 107.280 69.640 107.540 ;
        RECT 66.425 107.040 66.785 107.280 ;
        RECT 69.280 107.040 69.640 107.280 ;
        RECT 71.250 107.235 71.850 108.695 ;
        RECT 74.920 107.895 75.580 108.280 ;
        RECT 72.625 107.635 75.580 107.895 ;
        RECT 71.240 106.975 71.850 107.235 ;
        RECT 65.220 106.335 66.320 106.615 ;
        RECT 67.555 106.250 67.915 106.490 ;
        RECT 67.555 105.990 69.640 106.250 ;
        RECT 69.280 105.330 69.640 105.990 ;
        RECT 68.280 104.960 68.640 105.200 ;
        RECT 64.095 104.410 64.700 104.670 ;
        RECT 66.425 104.700 68.640 104.960 ;
        RECT 66.425 104.460 66.785 104.700 ;
        RECT 60.215 103.765 63.440 104.025 ;
        RECT 60.215 96.280 61.185 103.765 ;
        RECT 64.100 103.360 64.700 104.410 ;
        RECT 69.745 103.735 70.845 104.055 ;
        RECT 64.085 103.100 64.700 103.360 ;
        RECT 62.340 99.865 63.440 100.185 ;
        RECT 64.100 96.905 64.700 103.100 ;
        RECT 67.555 102.380 67.915 102.620 ;
        RECT 66.425 102.120 67.915 102.380 ;
        RECT 66.425 101.755 66.785 102.120 ;
        RECT 65.220 101.175 66.320 101.455 ;
        RECT 68.280 101.090 68.640 101.330 ;
        RECT 68.280 100.830 69.640 101.090 ;
        RECT 69.280 100.590 69.640 100.830 ;
        RECT 71.250 99.500 71.850 106.975 ;
        RECT 72.625 105.045 73.725 105.325 ;
        RECT 72.625 102.465 73.725 102.745 ;
        RECT 74.920 100.155 75.580 107.635 ;
        RECT 72.625 99.895 75.580 100.155 ;
        RECT 71.250 99.240 71.860 99.500 ;
        RECT 65.220 98.595 66.320 98.875 ;
        RECT 67.555 98.510 67.915 98.750 ;
        RECT 67.555 98.250 69.640 98.510 ;
        RECT 69.280 97.590 69.640 98.250 ;
        RECT 68.280 97.220 68.640 97.460 ;
        RECT 64.095 96.645 64.700 96.905 ;
        RECT 66.425 96.960 68.640 97.220 ;
        RECT 66.425 96.720 66.785 96.960 ;
        RECT 60.215 96.020 63.440 96.280 ;
        RECT 60.215 88.545 61.185 96.020 ;
        RECT 64.100 95.645 64.700 96.645 ;
        RECT 69.745 95.995 70.845 96.315 ;
        RECT 64.100 95.385 64.710 95.645 ;
        RECT 62.340 92.125 63.440 92.445 ;
        RECT 64.100 89.180 64.700 95.385 ;
        RECT 67.555 94.640 67.915 94.880 ;
        RECT 66.425 94.380 67.915 94.640 ;
        RECT 66.425 94.010 66.785 94.380 ;
        RECT 65.220 93.435 66.320 93.715 ;
        RECT 71.250 93.705 71.850 99.240 ;
        RECT 72.625 97.305 73.725 97.585 ;
        RECT 72.625 94.725 73.725 95.005 ;
        RECT 68.280 93.350 68.640 93.590 ;
        RECT 71.245 93.445 71.850 93.705 ;
        RECT 68.280 93.090 69.640 93.350 ;
        RECT 69.280 92.850 69.640 93.090 ;
        RECT 71.250 93.020 71.850 93.445 ;
        RECT 71.250 92.760 71.860 93.020 ;
        RECT 65.220 90.855 66.320 91.135 ;
        RECT 67.555 90.770 67.915 91.010 ;
        RECT 67.555 90.510 69.640 90.770 ;
        RECT 69.280 89.850 69.640 90.510 ;
        RECT 68.280 89.480 68.640 89.720 ;
        RECT 66.425 89.220 68.640 89.480 ;
        RECT 64.100 88.920 64.705 89.180 ;
        RECT 66.425 88.980 66.785 89.220 ;
        RECT 60.215 88.285 63.440 88.545 ;
        RECT 60.215 80.805 61.185 88.285 ;
        RECT 64.100 87.870 64.700 88.920 ;
        RECT 69.745 88.255 70.845 88.575 ;
        RECT 64.095 87.610 64.700 87.870 ;
        RECT 62.340 84.385 63.440 84.705 ;
        RECT 60.215 80.545 63.440 80.805 ;
        RECT 60.215 75.895 61.185 80.545 ;
        RECT 64.100 79.255 64.700 87.610 ;
        RECT 67.555 86.900 67.915 87.140 ;
        RECT 66.425 86.640 67.915 86.900 ;
        RECT 66.425 86.240 66.785 86.640 ;
        RECT 65.220 85.695 66.320 85.975 ;
        RECT 68.280 85.610 68.640 85.850 ;
        RECT 68.280 85.350 69.640 85.610 ;
        RECT 69.280 85.110 69.640 85.350 ;
        RECT 71.250 85.280 71.850 92.760 ;
        RECT 74.920 92.415 75.580 99.895 ;
        RECT 72.625 92.155 75.580 92.415 ;
        RECT 72.625 89.565 73.725 89.845 ;
        RECT 72.625 86.985 73.725 87.265 ;
        RECT 71.240 85.020 71.850 85.280 ;
        RECT 71.250 84.000 71.850 85.020 ;
        RECT 74.920 84.675 75.580 92.155 ;
        RECT 78.630 84.835 79.685 112.335 ;
        RECT 82.880 112.245 83.380 115.405 ;
        RECT 82.880 111.985 85.080 112.245 ;
        RECT 82.880 111.920 83.380 111.985 ;
        RECT 80.430 111.660 83.380 111.920 ;
        RECT 80.430 106.500 80.830 111.660 ;
        RECT 81.010 109.340 81.410 110.630 ;
        RECT 86.570 109.955 87.425 112.485 ;
        RECT 84.630 109.695 87.425 109.955 ;
        RECT 81.010 109.080 85.075 109.340 ;
        RECT 81.010 107.790 81.410 109.080 ;
        RECT 86.570 107.050 87.425 109.695 ;
        RECT 84.625 106.790 87.425 107.050 ;
        RECT 86.570 105.715 87.425 106.790 ;
        RECT 80.430 100.050 80.830 105.470 ;
        RECT 81.010 102.890 81.410 104.180 ;
        RECT 81.010 102.630 85.030 102.890 ;
        RECT 81.010 101.340 81.410 102.630 ;
        RECT 86.600 100.600 87.395 105.715 ;
        RECT 84.630 100.340 87.395 100.600 ;
        RECT 80.430 93.890 80.830 99.020 ;
        RECT 81.010 96.440 81.410 97.730 ;
        RECT 81.010 96.180 85.030 96.440 ;
        RECT 81.010 94.890 81.410 96.180 ;
        RECT 86.600 94.150 87.395 100.340 ;
        RECT 84.630 93.890 87.395 94.150 ;
        RECT 80.430 93.570 80.850 93.890 ;
        RECT 80.430 87.150 80.830 92.570 ;
        RECT 81.010 89.990 81.410 91.280 ;
        RECT 86.600 90.655 87.395 93.890 ;
        RECT 101.855 93.515 102.250 127.480 ;
        RECT 103.810 127.450 126.555 128.000 ;
        RECT 103.985 127.415 126.555 127.450 ;
        RECT 110.600 126.235 121.240 126.850 ;
        RECT 110.600 123.545 110.890 126.235 ;
        RECT 113.470 125.460 113.730 125.465 ;
        RECT 118.050 125.460 118.310 125.465 ;
        RECT 113.470 124.960 122.710 125.460 ;
        RECT 113.470 124.565 113.730 124.960 ;
        RECT 115.660 123.825 116.130 124.610 ;
        RECT 118.050 124.565 118.310 124.960 ;
        RECT 111.065 122.535 111.535 123.320 ;
        RECT 120.240 122.535 120.710 123.320 ;
        RECT 112.375 122.020 113.375 122.380 ;
        RECT 114.665 122.020 115.665 122.380 ;
        RECT 116.955 122.020 117.955 122.380 ;
        RECT 119.245 122.020 120.245 122.380 ;
        RECT 103.680 121.160 104.095 121.760 ;
        RECT 112.875 121.160 113.375 122.020 ;
        RECT 103.630 120.230 104.195 120.830 ;
        RECT 111.535 119.895 112.035 120.830 ;
        RECT 113.825 119.895 114.325 121.760 ;
        RECT 115.165 120.230 115.665 122.020 ;
        RECT 116.115 119.895 116.615 121.760 ;
        RECT 117.455 120.230 117.955 122.020 ;
        RECT 119.745 121.160 120.245 122.020 ;
        RECT 118.405 119.895 118.905 120.830 ;
        RECT 111.535 119.535 112.535 119.895 ;
        RECT 113.825 119.535 114.825 119.895 ;
        RECT 116.115 119.535 117.115 119.895 ;
        RECT 118.405 119.535 119.405 119.895 ;
        RECT 111.070 118.590 111.540 119.375 ;
        RECT 120.230 118.590 120.700 119.375 ;
        RECT 106.735 118.000 108.295 118.050 ;
        RECT 110.555 118.000 110.925 118.465 ;
        RECT 106.735 116.910 110.925 118.000 ;
        RECT 115.655 117.535 116.125 118.320 ;
        RECT 106.735 116.860 108.295 116.910 ;
        RECT 110.555 115.310 110.925 116.910 ;
        RECT 113.470 116.965 113.730 117.350 ;
        RECT 118.050 116.965 118.310 117.350 ;
        RECT 122.210 116.965 122.710 124.960 ;
        RECT 126.035 124.875 126.555 127.415 ;
        RECT 126.035 124.165 128.960 124.875 ;
        RECT 126.035 121.620 126.555 124.165 ;
        RECT 126.920 123.775 127.180 124.165 ;
        RECT 128.700 123.775 128.960 124.165 ;
        RECT 127.560 119.970 127.820 123.395 ;
        RECT 129.340 121.245 129.600 123.395 ;
        RECT 148.535 121.245 149.430 121.295 ;
        RECT 129.340 120.345 149.430 121.245 ;
        RECT 129.340 119.395 129.600 120.345 ;
        RECT 127.120 117.550 127.380 119.325 ;
        RECT 128.900 117.550 129.160 119.325 ;
        RECT 113.470 116.465 122.710 116.965 ;
        RECT 113.470 116.450 113.730 116.465 ;
        RECT 118.050 116.450 118.705 116.465 ;
        RECT 110.330 115.275 111.465 115.310 ;
        RECT 110.330 114.325 117.045 115.275 ;
        RECT 110.330 112.085 112.020 114.325 ;
        RECT 118.095 113.880 118.705 116.450 ;
        RECT 123.055 116.090 129.945 117.550 ;
        RECT 123.505 115.090 124.210 115.140 ;
        RECT 123.505 114.780 125.545 115.090 ;
        RECT 130.755 115.085 131.115 120.345 ;
        RECT 148.535 120.290 149.430 120.345 ;
        RECT 123.505 114.730 124.210 114.780 ;
        RECT 124.535 114.730 125.545 114.780 ;
        RECT 128.705 114.725 131.115 115.085 ;
        RECT 116.665 113.455 118.710 113.880 ;
        RECT 112.855 112.615 113.135 113.415 ;
        RECT 110.330 111.665 115.830 112.085 ;
        RECT 110.330 109.495 112.020 111.665 ;
        RECT 118.095 110.300 118.705 113.455 ;
        RECT 116.665 109.875 118.710 110.300 ;
        RECT 110.120 109.380 112.020 109.495 ;
        RECT 119.775 109.380 120.830 114.635 ;
        RECT 110.120 108.085 120.830 109.380 ;
        RECT 110.120 108.075 111.465 108.085 ;
        RECT 110.120 108.070 110.920 108.075 ;
        RECT 119.775 108.030 120.830 108.085 ;
        RECT 90.495 90.655 92.605 90.705 ;
        RECT 81.010 89.730 85.030 89.990 ;
        RECT 81.010 88.440 81.410 89.730 ;
        RECT 86.600 88.715 92.605 90.655 ;
        RECT 86.600 87.700 87.395 88.715 ;
        RECT 90.495 88.665 92.605 88.715 ;
        RECT 151.810 88.235 152.710 103.925 ;
        RECT 84.630 87.440 87.395 87.700 ;
        RECT 72.625 84.415 75.580 84.675 ;
        RECT 71.245 83.740 71.850 84.000 ;
        RECT 65.220 83.115 66.320 83.395 ;
        RECT 67.555 83.030 67.915 83.270 ;
        RECT 67.555 82.770 69.640 83.030 ;
        RECT 69.280 82.030 69.640 82.770 ;
        RECT 68.280 81.740 68.640 81.980 ;
        RECT 66.425 81.480 68.640 81.740 ;
        RECT 66.425 81.240 66.785 81.480 ;
        RECT 69.745 80.515 70.845 80.835 ;
        RECT 67.555 79.160 67.915 79.400 ;
        RECT 66.425 78.900 67.915 79.160 ;
        RECT 66.425 78.660 66.785 78.900 ;
        RECT 65.220 77.955 66.320 78.235 ;
        RECT 68.280 77.870 68.640 78.110 ;
        RECT 68.280 77.610 69.640 77.870 ;
        RECT 69.280 77.370 69.640 77.610 ;
        RECT 71.250 77.610 71.850 83.740 ;
        RECT 72.625 81.825 73.725 82.105 ;
        RECT 74.920 81.700 75.580 84.415 ;
        RECT 80.430 84.030 80.830 86.120 ;
        RECT 86.600 85.145 87.395 87.440 ;
        RECT 151.790 87.385 152.730 88.235 ;
        RECT 151.810 87.360 152.710 87.385 ;
        RECT 86.600 85.140 87.935 85.145 ;
        RECT 84.365 84.260 85.165 84.580 ;
        RECT 76.820 83.630 80.830 84.030 ;
        RECT 86.030 83.260 87.935 85.140 ;
        RECT 84.545 83.000 87.935 83.260 ;
        RECT 74.920 80.930 82.535 81.700 ;
        RECT 84.365 81.680 85.165 82.000 ;
        RECT 72.620 79.245 73.720 79.525 ;
        RECT 74.920 79.170 75.580 80.930 ;
        RECT 77.850 79.705 80.950 80.075 ;
        RECT 71.250 77.350 71.860 77.610 ;
        RECT 71.250 77.230 71.850 77.350 ;
        RECT 62.340 76.645 63.440 76.965 ;
        RECT 74.920 76.935 76.305 79.170 ;
        RECT 72.625 76.675 76.305 76.935 ;
        RECT 74.920 76.510 76.305 76.675 ;
        RECT 81.585 76.535 82.535 80.930 ;
        RECT 83.765 78.745 84.190 80.540 ;
        RECT 86.030 80.210 87.935 83.000 ;
        RECT 86.040 78.635 87.935 80.210 ;
        RECT 84.365 78.375 87.935 78.635 ;
        RECT 74.920 75.895 75.190 76.510 ;
        RECT 60.215 75.625 75.190 75.895 ;
        RECT 78.775 75.730 82.535 76.535 ;
        RECT 83.765 76.475 84.190 78.270 ;
        RECT 86.040 77.335 87.935 78.375 ;
        RECT 85.945 77.075 87.935 77.335 ;
        RECT 60.215 75.050 61.185 75.625 ;
        RECT 86.040 75.245 87.935 77.075 ;
        RECT 86.370 75.240 87.935 75.245 ;
        RECT 87.115 74.890 87.935 75.240 ;
        RECT 69.815 61.365 70.840 61.415 ;
        RECT 39.225 59.460 70.840 61.365 ;
        RECT 9.515 52.100 11.515 52.150 ;
        RECT 13.390 52.100 14.360 52.795 ;
        RECT 39.225 52.400 41.130 59.460 ;
        RECT 69.815 59.410 70.840 59.460 ;
        RECT 129.510 57.025 130.680 57.070 ;
        RECT 88.630 55.025 130.680 57.025 ;
        RECT 9.515 52.020 14.360 52.100 ;
        RECT 9.515 51.750 28.365 52.020 ;
        RECT 9.515 50.100 14.360 51.750 ;
        RECT 28.095 51.135 28.365 51.750 ;
        RECT 15.515 50.680 16.615 51.000 ;
        RECT 28.095 50.970 29.480 51.135 ;
        RECT 31.950 51.110 35.710 51.915 ;
        RECT 39.215 51.900 41.130 52.400 ;
        RECT 25.800 50.710 29.480 50.970 ;
        RECT 24.425 50.295 25.025 50.415 ;
        RECT 9.515 50.050 11.515 50.100 ;
        RECT 13.390 47.100 14.360 50.100 ;
        RECT 22.455 50.035 22.815 50.275 ;
        RECT 21.455 49.775 22.815 50.035 ;
        RECT 24.425 50.035 25.035 50.295 ;
        RECT 18.395 49.410 19.495 49.690 ;
        RECT 21.455 49.535 21.815 49.775 ;
        RECT 19.600 48.745 19.960 48.985 ;
        RECT 19.600 48.485 21.090 48.745 ;
        RECT 13.390 46.840 16.615 47.100 ;
        RECT 13.390 39.360 14.360 46.840 ;
        RECT 15.515 42.940 16.615 43.260 ;
        RECT 17.275 40.035 17.875 48.390 ;
        RECT 20.730 48.245 21.090 48.485 ;
        RECT 22.920 46.810 24.020 47.130 ;
        RECT 19.600 46.165 19.960 46.405 ;
        RECT 19.600 45.905 21.815 46.165 ;
        RECT 21.455 45.665 21.815 45.905 ;
        RECT 22.455 44.875 22.815 45.615 ;
        RECT 20.730 44.615 22.815 44.875 ;
        RECT 18.395 44.250 19.495 44.530 ;
        RECT 20.730 44.375 21.090 44.615 ;
        RECT 24.425 43.905 25.025 50.035 ;
        RECT 28.095 48.475 29.480 50.710 ;
        RECT 25.795 48.120 26.895 48.400 ;
        RECT 28.095 46.715 28.755 48.475 ;
        RECT 31.025 47.570 34.125 47.940 ;
        RECT 34.760 46.715 35.710 51.110 ;
        RECT 36.940 49.375 37.365 51.170 ;
        RECT 39.215 50.570 41.110 51.900 ;
        RECT 39.120 50.310 41.110 50.570 ;
        RECT 39.215 49.270 41.110 50.310 ;
        RECT 37.540 49.010 41.110 49.270 ;
        RECT 36.940 47.105 37.365 48.900 ;
        RECT 39.215 47.435 41.110 49.010 ;
        RECT 28.095 45.945 35.710 46.715 ;
        RECT 25.800 45.540 26.900 45.820 ;
        RECT 24.420 43.645 25.025 43.905 ;
        RECT 24.425 42.625 25.025 43.645 ;
        RECT 28.095 43.230 28.755 45.945 ;
        RECT 37.540 45.645 38.340 45.965 ;
        RECT 39.205 44.645 41.110 47.435 ;
        RECT 90.660 47.310 91.090 50.890 ;
        RECT 109.115 49.100 109.385 55.025 ;
        RECT 129.510 54.970 130.680 55.025 ;
        RECT 90.660 46.790 92.255 47.310 ;
        RECT 94.750 46.795 96.555 47.295 ;
        RECT 120.070 46.795 121.895 47.295 ;
        RECT 37.720 44.385 41.110 44.645 ;
        RECT 29.935 43.330 34.005 43.730 ;
        RECT 25.800 42.970 28.755 43.230 ;
        RECT 22.455 42.295 22.815 42.535 ;
        RECT 24.415 42.365 25.025 42.625 ;
        RECT 21.455 42.035 22.815 42.295 ;
        RECT 18.395 41.670 19.495 41.950 ;
        RECT 21.455 41.795 21.815 42.035 ;
        RECT 19.600 41.005 19.960 41.405 ;
        RECT 19.600 40.745 21.090 41.005 ;
        RECT 20.730 40.505 21.090 40.745 ;
        RECT 17.270 39.775 17.875 40.035 ;
        RECT 13.390 39.100 16.615 39.360 ;
        RECT 13.390 31.625 14.360 39.100 ;
        RECT 17.275 38.725 17.875 39.775 ;
        RECT 22.920 39.070 24.020 39.390 ;
        RECT 17.275 38.465 17.880 38.725 ;
        RECT 15.515 35.200 16.615 35.520 ;
        RECT 17.275 32.260 17.875 38.465 ;
        RECT 19.600 38.425 19.960 38.665 ;
        RECT 19.600 38.165 21.815 38.425 ;
        RECT 21.455 37.925 21.815 38.165 ;
        RECT 22.455 37.135 22.815 37.795 ;
        RECT 20.730 36.875 22.815 37.135 ;
        RECT 18.395 36.510 19.495 36.790 ;
        RECT 20.730 36.635 21.090 36.875 ;
        RECT 24.425 34.885 25.025 42.365 ;
        RECT 25.800 40.380 26.900 40.660 ;
        RECT 25.800 37.800 26.900 38.080 ;
        RECT 28.095 35.490 28.755 42.970 ;
        RECT 25.800 35.230 28.755 35.490 ;
        RECT 22.455 34.555 22.815 34.795 ;
        RECT 21.455 34.295 22.815 34.555 ;
        RECT 24.425 34.625 25.035 34.885 ;
        RECT 18.395 33.930 19.495 34.210 ;
        RECT 21.455 34.055 21.815 34.295 ;
        RECT 24.425 34.200 25.025 34.625 ;
        RECT 24.420 33.940 25.025 34.200 ;
        RECT 19.600 33.265 19.960 33.635 ;
        RECT 19.600 33.005 21.090 33.265 ;
        RECT 20.730 32.765 21.090 33.005 ;
        RECT 17.275 32.000 17.885 32.260 ;
        RECT 13.390 31.365 16.615 31.625 ;
        RECT 13.390 23.880 14.360 31.365 ;
        RECT 17.275 31.000 17.875 32.000 ;
        RECT 22.920 31.330 24.020 31.650 ;
        RECT 17.270 30.740 17.875 31.000 ;
        RECT 15.515 27.460 16.615 27.780 ;
        RECT 17.275 24.545 17.875 30.740 ;
        RECT 19.600 30.685 19.960 30.925 ;
        RECT 19.600 30.425 21.815 30.685 ;
        RECT 21.455 30.185 21.815 30.425 ;
        RECT 22.455 29.395 22.815 30.055 ;
        RECT 20.730 29.135 22.815 29.395 ;
        RECT 18.395 28.770 19.495 29.050 ;
        RECT 20.730 28.895 21.090 29.135 ;
        RECT 24.425 28.405 25.025 33.940 ;
        RECT 25.800 32.640 26.900 32.920 ;
        RECT 25.800 30.060 26.900 30.340 ;
        RECT 24.425 28.145 25.035 28.405 ;
        RECT 22.455 26.815 22.815 27.055 ;
        RECT 21.455 26.555 22.815 26.815 ;
        RECT 18.395 26.190 19.495 26.470 ;
        RECT 21.455 26.315 21.815 26.555 ;
        RECT 19.600 25.525 19.960 25.890 ;
        RECT 19.600 25.265 21.090 25.525 ;
        RECT 20.730 25.025 21.090 25.265 ;
        RECT 17.260 24.285 17.875 24.545 ;
        RECT 13.390 23.620 16.615 23.880 ;
        RECT 13.390 19.145 14.360 23.620 ;
        RECT 17.275 23.235 17.875 24.285 ;
        RECT 22.920 23.590 24.020 23.910 ;
        RECT 17.270 22.975 17.875 23.235 ;
        RECT 15.515 19.720 16.615 20.040 ;
        RECT 17.275 18.950 17.875 22.975 ;
        RECT 19.600 22.945 19.960 23.185 ;
        RECT 19.600 22.685 21.815 22.945 ;
        RECT 21.455 22.445 21.815 22.685 ;
        RECT 22.455 21.655 22.815 22.315 ;
        RECT 20.730 21.395 22.815 21.655 ;
        RECT 18.395 21.030 19.495 21.310 ;
        RECT 20.730 21.155 21.090 21.395 ;
        RECT 24.425 20.670 25.025 28.145 ;
        RECT 28.095 27.750 28.755 35.230 ;
        RECT 25.800 27.490 28.755 27.750 ;
        RECT 25.800 24.900 26.900 25.180 ;
        RECT 25.800 22.320 26.900 22.600 ;
        RECT 19.600 20.365 19.960 20.605 ;
        RECT 22.455 20.365 22.815 20.605 ;
        RECT 24.415 20.410 25.025 20.670 ;
        RECT 19.600 20.105 21.090 20.365 ;
        RECT 20.730 19.865 21.090 20.105 ;
        RECT 21.455 20.105 22.815 20.365 ;
        RECT 21.455 19.865 21.815 20.105 ;
        RECT 24.425 18.950 25.025 20.410 ;
        RECT 28.095 20.010 28.755 27.490 ;
        RECT 25.800 19.750 28.755 20.010 ;
        RECT 28.095 19.365 28.755 19.750 ;
        RECT 17.275 18.350 25.025 18.950 ;
        RECT 31.805 14.815 32.860 42.315 ;
        RECT 33.605 41.030 34.005 43.330 ;
        RECT 37.540 43.065 38.340 43.385 ;
        RECT 39.205 42.505 41.110 44.385 ;
        RECT 39.770 42.500 41.110 42.505 ;
        RECT 39.770 40.210 40.575 42.500 ;
        RECT 33.605 34.580 34.005 40.000 ;
        RECT 39.775 39.710 40.570 40.210 ;
        RECT 37.805 39.450 40.570 39.710 ;
        RECT 34.185 37.420 34.585 38.710 ;
        RECT 34.185 37.160 38.205 37.420 ;
        RECT 34.185 35.870 34.585 37.160 ;
        RECT 33.605 28.130 34.005 33.550 ;
        RECT 39.775 33.260 40.570 39.450 ;
        RECT 90.290 36.105 93.170 36.530 ;
        RECT 93.380 35.235 93.640 35.240 ;
        RECT 37.805 33.000 40.570 33.260 ;
        RECT 34.185 30.970 34.585 32.260 ;
        RECT 34.185 30.710 38.205 30.970 ;
        RECT 34.185 29.420 34.585 30.710 ;
        RECT 33.605 21.680 34.005 27.100 ;
        RECT 39.775 26.810 40.570 33.000 ;
        RECT 37.805 26.550 40.570 26.810 ;
        RECT 57.505 28.660 59.430 32.815 ;
        RECT 93.365 31.145 93.655 35.235 ;
        RECT 96.125 34.585 96.555 46.795 ;
        RECT 96.705 45.870 98.635 46.370 ;
        RECT 96.705 41.020 97.135 45.870 ;
        RECT 121.465 41.020 121.895 46.795 ;
        RECT 127.415 46.370 127.845 50.890 ;
        RECT 132.490 46.440 133.390 47.345 ;
        RECT 122.045 45.870 123.915 46.370 ;
        RECT 125.740 45.870 127.845 46.370 ;
        RECT 109.155 38.090 109.435 39.900 ;
        RECT 97.255 36.915 98.305 37.890 ;
        RECT 108.020 34.680 109.070 35.725 ;
        RECT 109.520 34.675 110.570 37.330 ;
        RECT 120.315 35.350 121.365 37.890 ;
        RECT 122.045 34.585 122.475 45.870 ;
        RECT 151.810 40.385 152.710 65.190 ;
        RECT 96.125 31.715 97.130 34.585 ;
        RECT 109.150 32.685 109.440 34.480 ;
        RECT 96.125 28.830 97.140 31.715 ;
        RECT 121.455 29.125 122.475 34.585 ;
        RECT 88.620 28.660 92.530 28.665 ;
        RECT 57.505 27.210 92.530 28.660 ;
        RECT 97.230 28.115 99.630 28.505 ;
        RECT 109.520 28.125 111.920 28.515 ;
        RECT 57.505 26.735 123.840 27.210 ;
        RECT 87.235 26.665 123.840 26.735 ;
        RECT 87.235 26.660 88.635 26.665 ;
        RECT 34.185 24.520 34.585 25.810 ;
        RECT 34.185 24.260 38.205 24.520 ;
        RECT 34.185 22.970 34.585 24.260 ;
        RECT 39.775 21.435 40.570 26.550 ;
        RECT 33.605 15.490 34.005 20.650 ;
        RECT 39.745 20.360 40.600 21.435 ;
        RECT 37.800 20.100 40.600 20.360 ;
        RECT 34.185 18.070 34.585 19.360 ;
        RECT 34.185 17.810 38.250 18.070 ;
        RECT 34.185 16.520 34.585 17.810 ;
        RECT 39.745 17.455 40.600 20.100 ;
        RECT 37.805 17.195 40.600 17.455 ;
        RECT 33.605 15.230 36.790 15.490 ;
        RECT 35.890 15.165 36.790 15.230 ;
        RECT 35.890 14.905 38.255 15.165 ;
        RECT 35.890 13.240 36.790 14.905 ;
        RECT 39.745 14.665 40.600 17.195 ;
      LAYER met3 ;
        RECT 59.275 164.355 71.770 164.940 ;
        RECT 54.625 154.780 58.375 155.630 ;
        RECT 64.945 154.315 65.365 158.910 ;
        RECT 64.945 153.860 70.905 154.315 ;
        RECT 65.015 153.815 70.905 153.860 ;
        RECT 60.560 147.675 60.980 152.725 ;
        RECT 69.325 147.675 69.745 152.725 ;
        RECT 70.405 142.735 70.905 153.815 ;
        RECT 82.820 149.735 93.220 156.490 ;
        RECT 82.820 148.835 133.070 149.735 ;
        RECT 82.820 146.250 93.220 148.835 ;
        RECT 76.595 145.700 93.220 146.250 ;
        RECT 82.820 144.630 93.220 145.700 ;
        RECT 70.405 142.720 71.360 142.735 ;
        RECT 60.565 142.220 71.360 142.720 ;
        RECT 36.555 135.435 36.945 138.805 ;
        RECT 60.565 137.670 60.985 142.220 ;
        RECT 69.325 137.670 69.745 142.220 ;
        RECT 17.695 135.060 36.945 135.435 ;
        RECT 15.025 125.570 15.615 127.620 ;
        RECT 20.770 125.295 21.670 134.140 ;
        RECT 36.555 131.640 36.945 135.060 ;
        RECT 64.945 131.870 65.365 136.920 ;
        RECT 24.635 127.070 27.135 127.410 ;
        RECT 36.925 127.080 39.425 127.420 ;
        RECT 20.720 124.775 21.720 125.295 ;
        RECT 20.770 124.300 21.670 124.775 ;
        RECT 24.635 64.850 25.535 127.070 ;
        RECT 36.925 68.925 37.825 127.080 ;
        RECT 60.580 122.040 61.070 122.590 ;
        RECT 70.810 121.710 71.360 142.220 ;
        RECT 115.755 136.625 116.175 137.675 ;
        RECT 105.175 135.745 105.595 136.295 ;
        RECT 126.335 135.745 126.755 136.295 ;
        RECT 105.175 135.245 128.955 135.745 ;
        RECT 105.175 130.815 105.595 131.865 ;
        RECT 126.335 130.815 126.755 131.865 ;
        RECT 115.755 129.935 116.175 130.485 ;
        RECT 128.455 129.935 128.955 135.245 ;
        RECT 115.755 129.435 128.955 129.935 ;
        RECT 115.610 123.850 116.180 124.585 ;
        RECT 121.605 123.295 122.340 129.435 ;
        RECT 99.235 122.040 99.875 122.590 ;
        RECT 111.015 122.560 122.340 123.295 ;
        RECT 103.630 121.710 104.145 121.735 ;
        RECT 70.810 121.160 101.725 121.710 ;
        RECT 103.475 121.210 104.145 121.710 ;
        RECT 103.630 121.185 104.145 121.210 ;
        RECT 101.175 120.780 101.725 121.160 ;
        RECT 103.580 120.780 104.245 120.805 ;
        RECT 79.915 119.990 80.490 120.540 ;
        RECT 101.175 120.280 104.245 120.780 ;
        RECT 101.175 119.660 101.725 120.280 ;
        RECT 103.580 120.255 104.245 120.280 ;
        RECT 60.615 119.110 101.725 119.660 ;
        RECT 111.020 118.615 111.590 119.350 ;
        RECT 120.180 118.615 120.750 119.350 ;
        RECT 115.605 118.270 116.175 118.295 ;
        RECT 121.605 118.270 122.340 122.560 ;
        RECT 45.595 116.885 46.965 118.025 ;
        RECT 59.300 116.930 96.675 117.995 ;
        RECT 99.245 116.885 100.265 118.020 ;
        RECT 106.685 116.885 108.345 118.025 ;
        RECT 115.605 117.560 122.340 118.270 ;
        RECT 82.830 114.430 83.430 115.380 ;
        RECT 123.455 114.755 124.260 115.115 ;
        RECT 82.830 113.390 83.430 113.415 ;
        RECT 82.830 112.890 113.185 113.390 ;
        RECT 82.830 112.865 83.430 112.890 ;
        RECT 112.805 112.640 113.185 112.890 ;
        RECT 132.170 112.160 133.070 148.835 ;
        RECT 135.090 138.895 136.680 140.880 ;
        RECT 148.485 120.315 149.480 121.270 ;
        RECT 62.365 107.555 63.415 107.975 ;
        RECT 122.015 107.295 140.875 112.160 ;
        RECT 120.905 106.760 140.875 107.295 ;
        RECT 57.580 104.815 58.465 106.730 ;
        RECT 65.245 106.285 66.295 106.665 ;
        RECT 65.915 105.965 66.295 106.285 ;
        RECT 65.915 101.505 66.285 105.965 ;
        RECT 72.650 104.995 73.700 105.375 ;
        RECT 69.770 103.685 70.820 104.105 ;
        RECT 73.320 102.795 73.700 104.995 ;
        RECT 72.650 102.415 73.700 102.795 ;
        RECT 65.245 101.125 66.295 101.505 ;
        RECT 62.365 99.815 63.415 100.235 ;
        RECT 65.915 98.925 66.285 101.125 ;
        RECT 65.245 98.545 66.295 98.925 ;
        RECT 65.915 93.765 66.285 98.545 ;
        RECT 73.320 97.635 73.700 102.415 ;
        RECT 72.650 97.255 73.700 97.635 ;
        RECT 69.770 95.945 70.820 96.365 ;
        RECT 73.320 95.055 73.700 97.255 ;
        RECT 72.650 94.675 73.700 95.055 ;
        RECT 122.015 94.760 140.875 106.760 ;
        RECT 151.760 103.135 152.760 103.900 ;
        RECT 65.245 93.385 66.295 93.765 ;
        RECT 62.365 92.075 63.415 92.495 ;
        RECT 65.915 91.185 66.285 93.385 ;
        RECT 65.245 90.805 66.295 91.185 ;
        RECT 65.915 86.025 66.285 90.805 ;
        RECT 73.320 89.895 73.700 94.675 ;
        RECT 80.455 93.520 81.040 93.940 ;
        RECT 101.720 93.510 102.335 93.930 ;
        RECT 72.650 89.515 73.700 89.895 ;
        RECT 69.770 88.205 70.820 88.625 ;
        RECT 73.320 87.315 73.700 89.515 ;
        RECT 90.445 88.690 92.655 90.680 ;
        RECT 151.815 88.260 152.705 88.285 ;
        RECT 151.810 87.360 152.710 88.260 ;
        RECT 151.815 87.335 152.705 87.360 ;
        RECT 72.650 86.935 73.700 87.315 ;
        RECT 65.245 85.645 66.295 86.025 ;
        RECT 62.365 84.335 63.415 84.755 ;
        RECT 65.915 83.445 66.285 85.645 ;
        RECT 65.245 83.065 66.295 83.445 ;
        RECT 65.915 78.285 66.285 83.065 ;
        RECT 73.320 82.535 73.700 86.935 ;
        RECT 84.390 84.210 85.140 84.630 ;
        RECT 76.845 83.580 77.260 84.080 ;
        RECT 76.870 82.535 77.235 83.580 ;
        RECT 73.320 82.155 77.235 82.535 ;
        RECT 72.650 81.775 73.700 82.155 ;
        RECT 69.770 80.465 70.820 80.885 ;
        RECT 73.320 79.575 73.700 81.775 ;
        RECT 84.390 81.630 85.140 82.050 ;
        RECT 77.875 79.655 80.925 80.125 ;
        RECT 72.645 79.195 73.700 79.575 ;
        RECT 65.245 77.905 66.295 78.285 ;
        RECT 62.365 76.595 63.415 77.015 ;
        RECT 65.915 76.325 66.285 77.905 ;
        RECT 73.320 76.325 73.700 79.195 ;
        RECT 83.790 78.695 84.165 80.590 ;
        RECT 83.790 76.425 84.165 78.320 ;
        RECT 65.915 75.955 73.700 76.325 ;
        RECT 36.925 68.025 58.910 68.925 ;
        RECT 24.635 63.950 47.135 64.850 ;
        RECT 151.760 64.430 152.760 65.165 ;
        RECT 69.765 59.435 70.890 61.390 ;
        RECT 24.335 55.870 59.430 57.795 ;
        RECT 9.465 50.075 11.565 52.125 ;
        RECT 19.090 51.320 26.875 51.690 ;
        RECT 15.540 50.630 16.590 51.050 ;
        RECT 19.090 49.740 19.460 51.320 ;
        RECT 18.420 49.360 19.470 49.740 ;
        RECT 19.090 44.580 19.460 49.360 ;
        RECT 26.495 48.450 26.875 51.320 ;
        RECT 36.965 49.325 37.340 51.220 ;
        RECT 25.820 48.070 26.875 48.450 ;
        RECT 22.945 46.760 23.995 47.180 ;
        RECT 26.495 45.870 26.875 48.070 ;
        RECT 31.050 47.520 34.100 47.990 ;
        RECT 36.965 47.055 37.340 48.950 ;
        RECT 25.825 45.490 26.875 45.870 ;
        RECT 37.565 45.595 38.315 46.015 ;
        RECT 26.495 45.110 30.410 45.490 ;
        RECT 18.420 44.200 19.470 44.580 ;
        RECT 15.540 42.890 16.590 43.310 ;
        RECT 19.090 42.000 19.460 44.200 ;
        RECT 18.420 41.620 19.470 42.000 ;
        RECT 19.090 36.840 19.460 41.620 ;
        RECT 26.495 40.710 26.875 45.110 ;
        RECT 29.985 43.780 30.410 45.110 ;
        RECT 29.960 43.280 30.435 43.780 ;
        RECT 37.565 43.015 38.315 43.435 ;
        RECT 25.825 40.330 26.875 40.710 ;
        RECT 22.945 39.020 23.995 39.440 ;
        RECT 26.495 38.130 26.875 40.330 ;
        RECT 25.825 37.750 26.875 38.130 ;
        RECT 18.420 36.460 19.470 36.840 ;
        RECT 15.540 35.150 16.590 35.570 ;
        RECT 19.090 34.260 19.460 36.460 ;
        RECT 18.420 33.880 19.470 34.260 ;
        RECT 19.090 29.100 19.460 33.880 ;
        RECT 26.495 32.970 26.875 37.750 ;
        RECT 25.825 32.590 26.875 32.970 ;
        RECT 57.505 32.795 59.430 55.870 ;
        RECT 129.460 54.995 130.730 57.045 ;
        RECT 132.440 46.490 133.440 47.315 ;
        RECT 151.760 40.410 152.760 41.175 ;
        RECT 109.100 36.505 109.490 39.875 ;
        RECT 90.240 36.130 109.490 36.505 ;
        RECT 22.945 31.280 23.995 31.700 ;
        RECT 26.495 30.390 26.875 32.590 ;
        RECT 57.480 30.820 59.455 32.795 ;
        RECT 25.825 30.010 26.875 30.390 ;
        RECT 18.420 28.720 19.470 29.100 ;
        RECT 15.540 27.410 16.590 27.830 ;
        RECT 19.090 26.520 19.460 28.720 ;
        RECT 18.420 26.140 19.470 26.520 ;
        RECT 19.090 21.680 19.460 26.140 ;
        RECT 26.495 25.230 26.875 30.010 ;
        RECT 25.825 24.850 26.875 25.230 ;
        RECT 22.945 23.540 23.995 23.960 ;
        RECT 26.495 22.650 26.875 24.850 ;
        RECT 25.825 22.270 26.875 22.650 ;
        RECT 19.090 21.360 19.470 21.680 ;
        RECT 18.420 20.980 19.470 21.360 ;
        RECT 15.540 19.670 16.590 20.090 ;
        RECT 93.315 17.855 94.215 35.210 ;
        RECT 109.100 32.710 109.490 36.130 ;
        RECT 74.530 16.955 94.215 17.855 ;
        RECT 97.180 28.140 99.680 28.480 ;
        RECT 109.470 28.150 111.970 28.490 ;
        RECT 35.840 13.265 36.840 13.860 ;
        RECT 74.530 9.090 75.430 16.955 ;
        RECT 97.180 14.025 98.080 28.140 ;
        RECT 109.470 21.505 110.370 28.150 ;
        RECT 109.420 20.605 110.420 21.505 ;
        RECT 109.470 20.595 110.370 20.605 ;
        RECT 97.130 13.125 98.130 14.025 ;
        RECT 74.480 8.190 75.480 9.090 ;
      LAYER met4 ;
        RECT 30.670 219.595 30.970 224.760 ;
        RECT 33.430 219.595 33.730 224.760 ;
        RECT 36.190 219.595 36.490 224.760 ;
        RECT 38.950 219.595 39.250 224.760 ;
        RECT 41.710 219.595 42.010 224.760 ;
        RECT 44.470 219.595 44.770 224.760 ;
        RECT 47.230 219.595 47.530 224.760 ;
        RECT 49.990 219.595 50.290 224.760 ;
        RECT 52.750 219.595 53.050 224.760 ;
        RECT 55.510 219.595 55.810 224.760 ;
        RECT 58.270 219.595 58.570 224.760 ;
        RECT 61.030 219.595 61.330 224.760 ;
        RECT 63.790 219.595 64.090 224.760 ;
        RECT 66.550 219.595 66.850 224.760 ;
        RECT 69.310 219.595 69.610 224.760 ;
        RECT 72.070 219.595 72.370 224.760 ;
        RECT 74.830 219.595 75.130 224.760 ;
        RECT 77.590 219.595 77.890 224.760 ;
        RECT 80.350 219.595 80.650 224.760 ;
        RECT 83.110 219.595 83.410 224.760 ;
        RECT 85.870 219.595 86.170 224.760 ;
        RECT 88.630 219.595 88.930 224.760 ;
        RECT 91.390 219.595 91.690 224.760 ;
        RECT 94.150 219.595 94.450 224.760 ;
        RECT 4.000 216.410 95.080 219.595 ;
        RECT 157.000 165.995 157.005 220.760 ;
        RECT 71.720 165.990 157.005 165.995 ;
        RECT 58.555 165.985 157.005 165.990 ;
        RECT 57.350 163.990 157.005 165.985 ;
        RECT 57.350 155.610 59.650 163.990 ;
        RECT 72.510 163.985 157.005 163.990 ;
        RECT 82.880 155.990 93.160 156.470 ;
        RECT 54.670 154.800 59.650 155.610 ;
        RECT 57.350 153.970 59.650 154.800 ;
        RECT 60.605 148.195 60.935 152.705 ;
        RECT 69.370 148.195 69.700 152.705 ;
        RECT 60.605 147.695 72.875 148.195 ;
        RECT 64.990 136.725 65.320 136.900 ;
        RECT 72.375 136.725 72.875 147.695 ;
        RECT 83.215 145.550 92.825 154.635 ;
        RECT 157.000 152.800 157.005 163.985 ;
        RECT 156.995 150.800 157.005 152.800 ;
        RECT 83.215 145.220 99.835 145.550 ;
        RECT 83.215 145.025 92.825 145.220 ;
        RECT 64.990 136.225 72.875 136.725 ;
        RECT 99.505 136.655 99.835 145.220 ;
        RECT 157.000 140.875 157.005 150.800 ;
        RECT 135.135 140.855 136.635 140.860 ;
        RECT 145.230 140.855 157.005 140.875 ;
        RECT 133.825 138.920 157.005 140.855 ;
        RECT 135.135 138.915 136.635 138.920 ;
        RECT 144.435 138.105 157.005 138.920 ;
        RECT 64.990 131.890 65.320 136.225 ;
        RECT 15.070 127.595 15.570 127.600 ;
        RECT 4.000 125.595 15.945 127.595 ;
        RECT 15.070 125.590 15.570 125.595 ;
        RECT 20.765 124.770 21.675 125.300 ;
        RECT 20.770 124.185 21.670 124.770 ;
        RECT 20.770 123.285 51.440 124.185 ;
        RECT 45.640 118.000 46.920 118.005 ;
        RECT 4.000 116.910 46.920 118.000 ;
        RECT 40.785 106.705 42.650 116.910 ;
        RECT 45.640 116.905 46.920 116.910 ;
        RECT 50.540 115.355 51.440 123.285 ;
        RECT 72.375 122.570 72.875 136.225 ;
        RECT 99.500 136.265 99.835 136.655 ;
        RECT 102.960 137.155 116.130 137.655 ;
        RECT 99.500 122.570 99.830 136.265 ;
        RECT 102.960 131.845 103.460 137.155 ;
        RECT 115.800 136.645 116.130 137.155 ;
        RECT 102.960 131.345 126.710 131.845 ;
        RECT 105.220 130.835 105.550 131.345 ;
        RECT 109.685 124.565 110.380 131.345 ;
        RECT 126.380 130.835 126.710 131.345 ;
        RECT 109.685 123.870 116.245 124.565 ;
        RECT 60.660 122.060 103.065 122.570 ;
        RECT 102.555 121.710 103.065 122.060 ;
        RECT 103.675 121.710 104.100 121.715 ;
        RECT 102.555 121.210 104.100 121.710 ;
        RECT 102.555 120.520 103.065 121.210 ;
        RECT 103.675 121.205 104.100 121.210 ;
        RECT 103.625 120.780 104.200 120.785 ;
        RECT 80.040 120.010 103.065 120.520 ;
        RECT 103.505 120.280 104.200 120.780 ;
        RECT 103.625 120.275 104.200 120.280 ;
        RECT 109.685 119.330 110.380 123.870 ;
        RECT 109.685 118.635 120.705 119.330 ;
        RECT 106.730 118.000 108.300 118.005 ;
        RECT 96.440 117.975 110.655 118.000 ;
        RECT 59.345 116.950 110.655 117.975 ;
        RECT 96.440 116.920 110.655 116.950 ;
        RECT 98.365 116.910 110.655 116.920 ;
        RECT 99.290 116.905 100.220 116.910 ;
        RECT 106.730 116.905 108.300 116.910 ;
        RECT 82.875 115.355 83.385 115.360 ;
        RECT 50.540 114.455 83.435 115.355 ;
        RECT 123.460 115.090 124.215 115.110 ;
        RECT 123.460 114.780 124.555 115.090 ;
        RECT 123.460 114.760 124.215 114.780 ;
        RECT 82.875 114.450 83.385 114.455 ;
        RECT 123.460 111.765 124.015 114.760 ;
        RECT 62.385 107.600 63.395 107.930 ;
        RECT 57.625 106.705 58.420 106.710 ;
        RECT 40.785 104.840 58.420 106.705 ;
        RECT 57.625 104.835 58.420 104.840 ;
        RECT 62.385 100.190 62.765 107.600 ;
        RECT 69.790 103.730 70.800 104.060 ;
        RECT 62.385 99.860 63.395 100.190 ;
        RECT 62.385 92.450 62.765 99.860 ;
        RECT 69.790 96.320 70.170 103.730 ;
        RECT 69.790 95.990 70.800 96.320 ;
        RECT 62.385 92.120 63.395 92.450 ;
        RECT 62.385 84.710 62.765 92.120 ;
        RECT 69.790 88.580 70.170 95.990 ;
        RECT 122.410 95.155 139.020 111.765 ;
        RECT 140.375 94.820 140.855 112.100 ;
        RECT 144.435 95.220 146.370 138.105 ;
        RECT 148.530 121.245 149.435 121.250 ;
        RECT 148.530 120.345 152.710 121.245 ;
        RECT 148.530 120.335 149.435 120.345 ;
        RECT 151.810 103.880 152.710 120.345 ;
        RECT 151.805 103.155 152.715 103.880 ;
        RECT 157.000 99.260 157.005 138.105 ;
        RECT 157.000 95.220 157.005 96.825 ;
        RECT 101.850 93.895 102.255 93.900 ;
        RECT 80.475 93.565 102.255 93.895 ;
        RECT 101.850 93.560 102.255 93.565 ;
        RECT 144.435 92.450 157.005 95.220 ;
        RECT 90.490 90.655 92.610 90.660 ;
        RECT 144.435 90.655 146.370 92.450 ;
        RECT 90.490 88.720 146.370 90.655 ;
        RECT 90.490 88.710 92.610 88.720 ;
        RECT 69.790 88.250 70.800 88.580 ;
        RECT 62.385 84.380 63.395 84.710 ;
        RECT 62.385 76.970 62.765 84.380 ;
        RECT 69.790 80.840 70.170 88.250 ;
        RECT 82.885 84.255 85.120 84.585 ;
        RECT 82.885 83.310 83.265 84.255 ;
        RECT 80.545 82.980 83.265 83.310 ;
        RECT 69.790 80.510 70.800 80.840 ;
        RECT 62.385 76.640 63.395 76.970 ;
        RECT 62.385 75.605 62.765 76.640 ;
        RECT 69.790 75.605 70.170 80.510 ;
        RECT 80.545 80.080 80.925 82.980 ;
        RECT 82.885 82.005 83.265 82.980 ;
        RECT 82.885 81.675 85.120 82.005 ;
        RECT 77.895 79.700 80.925 80.080 ;
        RECT 62.385 75.225 70.170 75.605 ;
        RECT 66.040 74.665 66.425 75.225 ;
        RECT 83.790 74.665 84.155 80.730 ;
        RECT 66.040 74.285 84.155 74.665 ;
        RECT 58.110 68.925 58.865 68.930 ;
        RECT 58.110 68.025 65.025 68.925 ;
        RECT 58.110 68.020 58.865 68.025 ;
        RECT 46.195 64.850 47.090 64.855 ;
        RECT 46.195 63.950 52.735 64.850 ;
        RECT 46.195 63.945 47.090 63.950 ;
        RECT 24.360 57.795 26.295 57.800 ;
        RECT 4.000 55.870 26.295 57.795 ;
        RECT 24.360 55.865 26.295 55.870 ;
        RECT 19.215 52.980 37.330 53.360 ;
        RECT 19.215 52.420 19.600 52.980 ;
        RECT 9.510 52.100 11.520 52.105 ;
        RECT 4.000 50.100 11.520 52.100 ;
        RECT 9.510 50.095 11.520 50.100 ;
        RECT 15.560 52.040 23.345 52.420 ;
        RECT 15.560 51.005 15.940 52.040 ;
        RECT 15.560 50.675 16.570 51.005 ;
        RECT 15.560 43.265 15.940 50.675 ;
        RECT 22.965 47.135 23.345 52.040 ;
        RECT 31.070 47.565 34.100 47.945 ;
        RECT 22.965 46.805 23.975 47.135 ;
        RECT 15.560 42.935 16.570 43.265 ;
        RECT 15.560 35.525 15.940 42.935 ;
        RECT 22.965 39.395 23.345 46.805 ;
        RECT 33.720 44.665 34.100 47.565 ;
        RECT 36.965 46.915 37.330 52.980 ;
        RECT 36.060 45.640 38.295 45.970 ;
        RECT 36.060 44.665 36.440 45.640 ;
        RECT 33.720 44.335 36.440 44.665 ;
        RECT 36.060 43.390 36.440 44.335 ;
        RECT 36.060 43.060 38.295 43.390 ;
        RECT 22.965 39.065 23.975 39.395 ;
        RECT 15.560 35.195 16.570 35.525 ;
        RECT 15.560 27.785 15.940 35.195 ;
        RECT 22.965 31.655 23.345 39.065 ;
        RECT 22.965 31.325 23.975 31.655 ;
        RECT 15.560 27.455 16.570 27.785 ;
        RECT 15.560 20.045 15.940 27.455 ;
        RECT 22.965 23.915 23.345 31.325 ;
        RECT 22.965 23.585 23.975 23.915 ;
        RECT 15.560 19.715 16.570 20.045 ;
        RECT 51.835 14.025 52.735 63.950 ;
        RECT 64.125 21.505 65.025 68.025 ;
        RECT 151.810 65.145 152.710 88.260 ;
        RECT 151.805 64.450 152.715 65.145 ;
        RECT 69.810 61.365 70.845 61.370 ;
        RECT 69.810 59.460 139.665 61.365 ;
        RECT 69.810 59.455 70.845 59.460 ;
        RECT 129.505 57.020 130.685 57.025 ;
        RECT 137.760 57.020 139.665 59.460 ;
        RECT 157.000 57.020 157.005 92.450 ;
        RECT 129.505 55.020 157.005 57.020 ;
        RECT 129.505 55.015 130.685 55.020 ;
        RECT 132.485 46.510 133.395 47.295 ;
        RECT 109.465 21.505 110.375 21.510 ;
        RECT 64.125 20.605 114.070 21.505 ;
        RECT 109.465 20.600 110.375 20.605 ;
        RECT 97.175 14.025 98.085 14.030 ;
        RECT 35.885 13.285 36.795 13.840 ;
        RECT 35.890 8.415 36.790 13.285 ;
        RECT 51.835 13.125 98.085 14.025 ;
        RECT 35.890 7.515 56.110 8.415 ;
        RECT 74.525 8.185 75.435 9.095 ;
        RECT 55.210 1.690 56.110 7.515 ;
        RECT 55.205 1.000 56.110 1.690 ;
        RECT 74.530 1.000 75.430 8.185 ;
        RECT 93.850 1.000 94.750 13.125 ;
        RECT 97.175 13.120 98.085 13.125 ;
        RECT 113.170 1.000 114.070 20.605 ;
        RECT 132.490 1.000 133.390 46.510 ;
        RECT 151.805 40.430 152.715 41.155 ;
        RECT 151.810 1.000 152.710 40.430 ;
        RECT 157.000 5.000 157.005 55.020 ;
        RECT 55.205 0.995 55.210 1.000 ;
  END
END tt_um_DalinEM_diff_amp
END LIBRARY

