magic
tech sky130A
magscale 1 2
timestamp 1741224942
<< metal1 >>
rect -2225 3760 -2001 3860
rect -2237 3451 -1997 3551
rect 7112 -1143 7122 -1043
rect 7205 -1143 7890 -1043
rect 7102 -1329 7112 -1229
rect 7225 -1329 7886 -1229
<< via1 >>
rect 7122 -1143 7205 -1043
rect 7112 -1329 7225 -1229
<< metal2 >>
rect -1749 7598 730 7608
rect -1749 7481 730 7491
rect -2376 5405 -1696 5808
rect 13414 2786 13712 2796
rect 5125 2443 7137 2786
rect 5125 2396 7293 2443
rect 12075 2399 13414 2785
rect 5125 2068 5524 2396
rect 7078 2368 7293 2396
rect 13414 2389 13712 2399
rect -10599 134 -10501 144
rect -10501 -266 -10349 134
rect -10599 -276 -10501 -266
rect -3764 -490 -3355 -167
rect -3767 -827 -1621 -490
rect 7122 -1043 7205 -1033
rect 7122 -1153 7205 -1143
rect 7112 -1229 7225 -1219
rect 12254 -1316 14187 -1136
rect 7112 -1339 7225 -1329
rect 6245 -1786 6429 -1776
rect 7733 -1785 8045 -1775
rect -1572 -3871 -1377 -1809
rect 6059 -2003 6245 -1786
rect 6429 -2003 6438 -1786
rect 6245 -2013 6429 -2003
rect 2962 -2314 3062 -2304
rect 2962 -2707 3062 -2494
rect 2962 -3053 3062 -2807
rect 6757 -6606 6836 -1934
rect 8045 -2003 8517 -1785
rect 7733 -2013 8045 -2003
rect 6757 -6682 6836 -6672
rect 4485 -7254 4907 -7244
rect 3786 -7642 4485 -7254
rect 4485 -7652 4907 -7642
<< via2 >>
rect -1749 7491 730 7598
rect 13414 2399 13712 2786
rect -10599 -266 -10501 134
rect 7122 -1143 7205 -1043
rect 7112 -1329 7225 -1229
rect 6245 -2003 6429 -1786
rect 2962 -2494 3062 -2314
rect 2962 -2807 3062 -2707
rect 7733 -2003 8045 -1785
rect 6757 -6672 6836 -6606
rect 4485 -7642 4907 -7254
<< metal3 >>
rect -1759 7598 740 7603
rect -1759 7491 -1749 7598
rect 730 7491 740 7598
rect -1759 7486 740 7491
rect 4941 4382 13000 4562
rect -10609 134 -10491 139
rect -10609 -266 -10599 134
rect -10501 -266 -10491 134
rect -10609 -271 -10491 -266
rect -9470 -430 -9460 -326
rect -9280 -430 -9270 -326
rect -9460 -525 -9280 -430
rect -8687 -991 -8507 -259
rect -6229 -958 -6049 -263
rect 7112 -1043 7215 -1038
rect 7081 -1143 7122 -1043
rect 7205 -1143 7215 -1043
rect 7112 -1148 7215 -1143
rect 7102 -1229 7235 -1224
rect 7102 -1329 7112 -1229
rect 7225 -1329 7235 -1229
rect 7102 -1334 7235 -1329
rect 6235 -1786 6439 -1781
rect 6235 -2003 6245 -1786
rect 6429 -2003 6439 -1786
rect 6235 -2008 6439 -2003
rect 7723 -1785 8055 -1780
rect 7723 -2003 7733 -1785
rect 8045 -2003 8055 -1785
rect 7723 -2008 8055 -2003
rect 2952 -2314 3072 -2309
rect 2952 -2494 2962 -2314
rect 3062 -2494 3072 -2314
rect 2952 -2499 3072 -2494
rect 2952 -2707 3072 -2702
rect 2952 -2807 2962 -2707
rect 3062 -2807 9013 -2707
rect 2952 -2812 3072 -2807
rect 12820 -3015 13000 4382
rect 13404 2786 13722 2791
rect 13404 2399 13414 2786
rect 13712 2399 13722 2786
rect 13404 2394 13722 2399
rect 6730 -6606 6853 -6599
rect 6730 -6672 6757 -6606
rect 6836 -6672 6853 -6606
rect 6730 -6683 6853 -6672
rect 4475 -7254 4917 -7249
rect 4475 -7642 4485 -7254
rect 4907 -7642 4917 -7254
rect 4475 -7647 4917 -7642
<< via3 >>
rect -1749 7491 730 7598
rect -10599 -266 -10501 134
rect -9460 -430 -9280 -326
rect 7122 -1143 7205 -1043
rect 7112 -1329 7225 -1229
rect 6245 -2003 6429 -1786
rect 7733 -2003 8045 -1785
rect 2962 -2494 3062 -2314
rect 13414 2399 13712 2786
rect 6757 -6672 6836 -6606
rect 4485 -7642 4907 -7254
<< metal4 >>
rect -1903 7598 897 7813
rect -1903 7491 -1749 7598
rect 730 7491 897 7598
rect -1903 7413 897 7491
rect 13413 2786 13713 2787
rect 13151 2399 13414 2786
rect 13712 2399 15660 2786
rect 13413 2398 13713 2399
rect -10600 134 -10500 135
rect -10693 -266 -10599 134
rect -10501 -266 -10425 134
rect -10600 -267 -10500 -266
rect -9461 -326 -9279 -325
rect -9461 -430 -9460 -326
rect -9280 -430 -9279 -326
rect -9461 -431 -9279 -430
rect -9460 -548 -9280 -431
rect -9460 -728 -3326 -548
rect -3506 -2314 -3326 -728
rect 7121 -1043 7206 -1042
rect 7121 -1143 7122 -1043
rect 7205 -1143 7206 -1043
rect 7121 -1144 7206 -1143
rect 7111 -1229 7226 -1228
rect 7087 -1329 7112 -1229
rect 7225 -1329 7226 -1229
rect 7111 -1330 7226 -1329
rect 7732 -1785 8046 -1784
rect 6244 -1786 7733 -1785
rect 6059 -2003 6245 -1786
rect 6429 -2003 7733 -1786
rect 8045 -2003 8517 -1785
rect 6244 -2004 6430 -2003
rect 7732 -2004 8046 -2003
rect 2961 -2314 3063 -2313
rect -3506 -2494 2962 -2314
rect 3062 -2494 3073 -2314
rect 2961 -2495 3063 -2494
rect 6756 -6606 6837 -6605
rect 4069 -6672 6757 -6606
rect 6836 -6672 6837 -6606
rect 6756 -6673 6837 -6672
rect 4484 -7254 4908 -7253
rect 15273 -7254 15660 2399
rect 4484 -7642 4485 -7254
rect 4907 -7641 15660 -7254
rect 4907 -7642 4908 -7641
rect 4484 -7643 4908 -7642
use 2nd_3_OTA  2nd_3_OTA_0 ~/Project_tinytape/magic/mag/OTA_stage2
timestamp 1741224555
transform 1 0 -8305 0 1 3126
box 6296 -5137 15454 4514
use 3rd_3_OTA  3rd_3_OTA_0 ~/Project_tinytape/magic/mag/3rd_3_OTA
timestamp 1741211560
transform 1 0 7949 0 -1 3001
box -1013 -144 6612 9434
use OTA_stage1  OTA_stage1_0 ~/Project_tinytape/magic/mag/OTA_stage1
timestamp 1741208255
transform 1 0 -21392 0 1 2425
box 10993 -2832 19171 3381
use OTA_vref  OTA_vref_0 ~/Project_tinytape/magic/mag/OTA_vref
timestamp 1740539468
transform 0 -1 4009 1 0 -10528
box 0 -73 7756 5648
<< labels >>
rlabel metal2 14185 -1227 14185 -1227 3 vo3
port 1 e
rlabel metal3 -6150 -956 -6150 -956 5 vin_p
port 2 s
rlabel metal3 -8592 -989 -8592 -989 5 vin_n
port 3 s
rlabel metal4 895 7673 895 7673 3 vcc
port 4 e
rlabel metal4 -10692 -78 -10692 -78 7 vss
port 5 w
<< end >>
