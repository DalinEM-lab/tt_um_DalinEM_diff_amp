magic
tech sky130A
magscale 1 2
timestamp 1741312032
<< nwell >>
rect 3323 29327 11333 30802
rect 11781 25249 14394 33008
rect 16817 25378 18823 27216
rect 20743 25468 25637 27902
rect 25243 24238 26061 25196
rect 16668 21223 17303 22596
rect 16652 19927 17290 20719
rect 16652 18637 17290 19429
rect 16652 17347 17290 18139
rect 16659 16222 17291 17053
rect 16658 15042 17291 16222
rect 16658 15038 17290 15042
rect 7293 10487 7925 10491
rect 7293 9307 7926 10487
rect 17832 9541 25842 11016
rect 7294 8476 7926 9307
rect 7287 7291 7925 8083
rect 7287 6001 7925 6793
rect 7287 4711 7925 5503
rect 7303 2834 7938 4207
<< pwell >>
rect 3327 25813 4347 27205
rect 4587 25282 10114 28837
rect 4671 25248 4694 25282
rect 4788 25248 10021 25250
rect 22119 23048 24255 25333
rect 12050 17216 15164 21866
rect 12050 17184 13294 17216
rect 13298 17215 15164 17216
rect 13298 17184 13344 17215
rect 12050 17182 13344 17184
rect 13347 17182 15164 17215
rect 12050 15024 15164 17182
rect 15760 16936 16607 22610
rect 22444 21850 23964 22900
rect 24723 22780 26127 23182
rect 15210 16265 16550 16418
rect 15210 15231 15363 16265
rect 16397 15231 16550 16265
rect 15210 15078 16550 15231
rect 2685 8347 5799 10505
rect 5845 10298 7185 10451
rect 5845 9264 5998 10298
rect 7032 9264 7185 10298
rect 5845 9111 7185 9264
rect 2685 8345 3979 8347
rect 2685 8313 3929 8345
rect 3933 8314 3979 8345
rect 3982 8314 5799 8347
rect 3933 8313 5799 8314
rect 2685 3663 5799 8313
rect 6395 2820 7242 8494
rect 17836 6027 18856 7419
rect 19096 5496 24623 9051
rect 19180 5462 19203 5496
rect 19297 5462 24530 5464
<< nbase >>
rect 15363 15231 16397 16265
rect 5998 9264 7032 10298
<< nmos >>
rect 3537 26009 4137 27009
rect 22654 22404 23754 22704
rect 22654 22046 23754 22346
rect 18046 6223 18646 7223
<< pmos >>
rect 17013 25597 17373 26997
rect 17431 25597 17791 26997
rect 17849 25597 18209 26997
rect 18267 25597 18627 26997
<< pmoslvt >>
rect 3712 30092 7312 30452
rect 7370 30092 10970 30452
rect 3712 29604 7312 29964
rect 7370 29604 10970 29964
rect 12184 29528 12564 32528
rect 12622 29528 13002 32528
rect 13060 29528 13440 32528
rect 13498 29528 13878 32528
rect 12184 25551 12564 28551
rect 12622 25551 13002 28551
rect 13060 25551 13440 28551
rect 13498 25551 13878 28551
rect 21106 27042 22106 27542
rect 22164 27042 23164 27542
rect 23222 27042 24222 27542
rect 24280 27042 25280 27542
rect 21106 25880 22106 26380
rect 22164 25880 23164 26380
rect 23222 25880 24222 26380
rect 24280 25880 25280 26380
rect 25439 24457 25509 24977
rect 25795 24457 25865 24977
rect 16871 21994 17071 22394
rect 16871 21413 17071 21813
rect 16871 20123 17071 20523
rect 16871 18833 17071 19233
rect 16871 17543 17071 17943
rect 16871 16655 17071 16855
rect 16871 16397 17071 16597
rect 16871 15730 16971 16130
rect 16871 15272 16971 15672
rect 7506 9857 7606 10257
rect 7506 9399 7606 9799
rect 7506 8932 7706 9132
rect 7506 8674 7706 8874
rect 18221 10306 21821 10666
rect 21879 10306 25479 10666
rect 18221 9818 21821 10178
rect 21879 9818 25479 10178
rect 7506 7487 7706 7887
rect 7506 6197 7706 6597
rect 7506 4907 7706 5307
rect 7506 3617 7706 4017
rect 7506 3036 7706 3436
<< nmoslvt >>
rect 4922 27380 7322 28580
rect 7380 27380 9780 28580
rect 4921 25505 7321 26705
rect 7379 25505 9779 26705
rect 12194 24225 14074 24525
rect 14132 24225 16012 24525
rect 16070 24225 17950 24525
rect 18008 24225 19888 24525
rect 12194 23815 14074 24115
rect 14132 23815 16012 24115
rect 16070 23815 17950 24115
rect 18008 23815 19888 24115
rect 22291 24495 22691 25095
rect 22749 24495 23149 25095
rect 23207 24495 23607 25095
rect 23665 24495 24065 25095
rect 22291 23288 22691 23888
rect 22749 23288 23149 23888
rect 23207 23288 23607 23888
rect 23665 23288 24065 23888
rect 25479 23772 25509 23972
rect 25835 23772 25865 23972
rect 12466 21324 13266 21524
rect 13947 21324 14747 21524
rect 12466 21066 13266 21266
rect 13947 21066 14747 21266
rect 12466 20808 13266 21008
rect 13947 20808 14747 21008
rect 12466 20550 13266 20750
rect 13947 20550 14747 20750
rect 12466 20292 13266 20492
rect 13947 20292 14747 20492
rect 12466 20034 13266 20234
rect 13947 20034 14747 20234
rect 12466 19776 13266 19976
rect 13947 19776 14747 19976
rect 12466 19518 13266 19718
rect 13947 19518 14747 19718
rect 12466 19260 13266 19460
rect 13947 19260 14747 19460
rect 12466 19002 13266 19202
rect 13947 19002 14747 19202
rect 12466 18744 13266 18944
rect 13947 18744 14747 18944
rect 12466 18486 13266 18686
rect 13947 18486 14747 18686
rect 12466 18228 13266 18428
rect 13947 18228 14747 18428
rect 12466 17970 13266 18170
rect 13947 17970 14747 18170
rect 12466 17712 13266 17912
rect 13947 17712 14747 17912
rect 12466 17454 13266 17654
rect 13947 17454 14747 17654
rect 12466 17196 13266 17396
rect 13947 17196 14747 17396
rect 12466 16938 13266 17138
rect 13947 16938 14747 17138
rect 12466 16680 13266 16880
rect 13947 16680 14747 16880
rect 12466 16422 13266 16622
rect 13947 16422 14747 16622
rect 12466 16164 13266 16364
rect 13947 16164 14747 16364
rect 12466 15906 13266 16106
rect 13947 15906 14747 16106
rect 12466 15648 13266 15848
rect 13947 15648 14747 15848
rect 12466 15390 13266 15590
rect 13947 15390 14747 15590
rect 16084 22129 16284 22329
rect 16084 21871 16284 22071
rect 16084 21613 16284 21813
rect 16084 21355 16284 21555
rect 16084 21097 16284 21297
rect 16084 20839 16284 21039
rect 16084 20581 16284 20781
rect 16084 20323 16284 20523
rect 16084 20065 16284 20265
rect 16084 19807 16284 20007
rect 16084 19549 16284 19749
rect 16084 19291 16284 19491
rect 16084 19033 16284 19233
rect 16084 18775 16284 18975
rect 16084 18517 16284 18717
rect 16084 18259 16284 18459
rect 16084 18001 16284 18201
rect 16084 17743 16284 17943
rect 16084 17485 16284 17685
rect 16084 17227 16284 17427
rect 3101 9939 3901 10139
rect 4582 9939 5382 10139
rect 3101 9681 3901 9881
rect 4582 9681 5382 9881
rect 3101 9423 3901 9623
rect 4582 9423 5382 9623
rect 3101 9165 3901 9365
rect 4582 9165 5382 9365
rect 3101 8907 3901 9107
rect 4582 8907 5382 9107
rect 3101 8649 3901 8849
rect 4582 8649 5382 8849
rect 3101 8391 3901 8591
rect 4582 8391 5382 8591
rect 3101 8133 3901 8333
rect 4582 8133 5382 8333
rect 3101 7875 3901 8075
rect 4582 7875 5382 8075
rect 3101 7617 3901 7817
rect 4582 7617 5382 7817
rect 3101 7359 3901 7559
rect 4582 7359 5382 7559
rect 3101 7101 3901 7301
rect 4582 7101 5382 7301
rect 3101 6843 3901 7043
rect 4582 6843 5382 7043
rect 3101 6585 3901 6785
rect 4582 6585 5382 6785
rect 3101 6327 3901 6527
rect 4582 6327 5382 6527
rect 3101 6069 3901 6269
rect 4582 6069 5382 6269
rect 3101 5811 3901 6011
rect 4582 5811 5382 6011
rect 3101 5553 3901 5753
rect 4582 5553 5382 5753
rect 3101 5295 3901 5495
rect 4582 5295 5382 5495
rect 3101 5037 3901 5237
rect 4582 5037 5382 5237
rect 3101 4779 3901 4979
rect 4582 4779 5382 4979
rect 3101 4521 3901 4721
rect 4582 4521 5382 4721
rect 3101 4263 3901 4463
rect 4582 4263 5382 4463
rect 3101 4005 3901 4205
rect 4582 4005 5382 4205
rect 6719 8003 6919 8203
rect 6719 7745 6919 7945
rect 6719 7487 6919 7687
rect 6719 7229 6919 7429
rect 6719 6971 6919 7171
rect 6719 6713 6919 6913
rect 6719 6455 6919 6655
rect 6719 6197 6919 6397
rect 6719 5939 6919 6139
rect 6719 5681 6919 5881
rect 6719 5423 6919 5623
rect 6719 5165 6919 5365
rect 6719 4907 6919 5107
rect 6719 4649 6919 4849
rect 6719 4391 6919 4591
rect 6719 4133 6919 4333
rect 6719 3875 6919 4075
rect 6719 3617 6919 3817
rect 6719 3359 6919 3559
rect 6719 3101 6919 3301
rect 19431 7594 21831 8794
rect 21889 7594 24289 8794
rect 19430 5719 21830 6919
rect 21888 5719 24288 6919
<< ndiff >>
rect 3537 27055 4137 27067
rect 3537 27021 3549 27055
rect 4125 27021 4137 27055
rect 3537 27009 4137 27021
rect 3537 25997 4137 26009
rect 3537 25963 3549 25997
rect 4125 25963 4137 25997
rect 3537 25951 4137 25963
rect 4864 28568 4922 28580
rect 4864 27392 4876 28568
rect 4910 27392 4922 28568
rect 4864 27380 4922 27392
rect 7322 28568 7380 28580
rect 7322 27392 7334 28568
rect 7368 27392 7380 28568
rect 7322 27380 7380 27392
rect 9780 28568 9838 28580
rect 9780 27392 9792 28568
rect 9826 27392 9838 28568
rect 9780 27380 9838 27392
rect 4863 26693 4921 26705
rect 4863 25517 4875 26693
rect 4909 25517 4921 26693
rect 4863 25505 4921 25517
rect 7321 26693 7379 26705
rect 7321 25517 7333 26693
rect 7367 25517 7379 26693
rect 7321 25505 7379 25517
rect 9779 26693 9837 26705
rect 9779 25517 9791 26693
rect 9825 25517 9837 26693
rect 9779 25505 9837 25517
rect 12136 24513 12194 24525
rect 12136 24237 12148 24513
rect 12182 24237 12194 24513
rect 12136 24225 12194 24237
rect 14074 24513 14132 24525
rect 14074 24237 14086 24513
rect 14120 24237 14132 24513
rect 14074 24225 14132 24237
rect 16012 24513 16070 24525
rect 16012 24237 16024 24513
rect 16058 24237 16070 24513
rect 16012 24225 16070 24237
rect 17950 24513 18008 24525
rect 17950 24237 17962 24513
rect 17996 24237 18008 24513
rect 17950 24225 18008 24237
rect 19888 24513 19946 24525
rect 19888 24237 19900 24513
rect 19934 24237 19946 24513
rect 19888 24225 19946 24237
rect 12136 24103 12194 24115
rect 12136 23827 12148 24103
rect 12182 23827 12194 24103
rect 12136 23815 12194 23827
rect 14074 24103 14132 24115
rect 14074 23827 14086 24103
rect 14120 23827 14132 24103
rect 14074 23815 14132 23827
rect 16012 24103 16070 24115
rect 16012 23827 16024 24103
rect 16058 23827 16070 24103
rect 16012 23815 16070 23827
rect 17950 24103 18008 24115
rect 17950 23827 17962 24103
rect 17996 23827 18008 24103
rect 17950 23815 18008 23827
rect 19888 24103 19946 24115
rect 19888 23827 19900 24103
rect 19934 23827 19946 24103
rect 19888 23815 19946 23827
rect 22233 25083 22291 25095
rect 22233 24507 22245 25083
rect 22279 24507 22291 25083
rect 22233 24495 22291 24507
rect 22691 25083 22749 25095
rect 22691 24507 22703 25083
rect 22737 24507 22749 25083
rect 22691 24495 22749 24507
rect 23149 25083 23207 25095
rect 23149 24507 23161 25083
rect 23195 24507 23207 25083
rect 23149 24495 23207 24507
rect 23607 25083 23665 25095
rect 23607 24507 23619 25083
rect 23653 24507 23665 25083
rect 23607 24495 23665 24507
rect 24065 25083 24123 25095
rect 24065 24507 24077 25083
rect 24111 24507 24123 25083
rect 24065 24495 24123 24507
rect 22233 23876 22291 23888
rect 22233 23300 22245 23876
rect 22279 23300 22291 23876
rect 22233 23288 22291 23300
rect 22691 23876 22749 23888
rect 22691 23300 22703 23876
rect 22737 23300 22749 23876
rect 22691 23288 22749 23300
rect 23149 23876 23207 23888
rect 23149 23300 23161 23876
rect 23195 23300 23207 23876
rect 23149 23288 23207 23300
rect 23607 23876 23665 23888
rect 23607 23300 23619 23876
rect 23653 23300 23665 23876
rect 23607 23288 23665 23300
rect 24065 23876 24123 23888
rect 24065 23300 24077 23876
rect 24111 23300 24123 23876
rect 24065 23288 24123 23300
rect 25421 23960 25479 23972
rect 25421 23784 25433 23960
rect 25467 23784 25479 23960
rect 25421 23772 25479 23784
rect 25509 23960 25567 23972
rect 25509 23784 25521 23960
rect 25555 23784 25567 23960
rect 25509 23772 25567 23784
rect 25777 23960 25835 23972
rect 25777 23784 25789 23960
rect 25823 23784 25835 23960
rect 25777 23772 25835 23784
rect 25865 23960 25923 23972
rect 25865 23784 25877 23960
rect 25911 23784 25923 23960
rect 25865 23772 25923 23784
rect 12466 21570 13266 21582
rect 12466 21536 12478 21570
rect 13254 21536 13266 21570
rect 12466 21524 13266 21536
rect 13947 21570 14747 21582
rect 13947 21536 13959 21570
rect 14735 21536 14747 21570
rect 13947 21524 14747 21536
rect 12466 21312 13266 21324
rect 12466 21278 12478 21312
rect 13254 21278 13266 21312
rect 12466 21266 13266 21278
rect 13947 21312 14747 21324
rect 13947 21278 13959 21312
rect 14735 21278 14747 21312
rect 13947 21266 14747 21278
rect 12466 21054 13266 21066
rect 12466 21020 12478 21054
rect 13254 21020 13266 21054
rect 12466 21008 13266 21020
rect 13947 21054 14747 21066
rect 13947 21020 13959 21054
rect 14735 21020 14747 21054
rect 13947 21008 14747 21020
rect 12466 20796 13266 20808
rect 12466 20762 12478 20796
rect 13254 20762 13266 20796
rect 12466 20750 13266 20762
rect 13947 20796 14747 20808
rect 13947 20762 13959 20796
rect 14735 20762 14747 20796
rect 13947 20750 14747 20762
rect 12466 20538 13266 20550
rect 12466 20504 12478 20538
rect 13254 20504 13266 20538
rect 12466 20492 13266 20504
rect 13947 20538 14747 20550
rect 13947 20504 13959 20538
rect 14735 20504 14747 20538
rect 13947 20492 14747 20504
rect 12466 20280 13266 20292
rect 12466 20246 12478 20280
rect 13254 20246 13266 20280
rect 12466 20234 13266 20246
rect 13947 20280 14747 20292
rect 13947 20246 13959 20280
rect 14735 20246 14747 20280
rect 13947 20234 14747 20246
rect 12466 20022 13266 20034
rect 12466 19988 12478 20022
rect 13254 19988 13266 20022
rect 12466 19976 13266 19988
rect 13947 20022 14747 20034
rect 13947 19988 13959 20022
rect 14735 19988 14747 20022
rect 13947 19976 14747 19988
rect 12466 19764 13266 19776
rect 12466 19730 12478 19764
rect 13254 19730 13266 19764
rect 12466 19718 13266 19730
rect 13947 19764 14747 19776
rect 13947 19730 13959 19764
rect 14735 19730 14747 19764
rect 13947 19718 14747 19730
rect 12466 19506 13266 19518
rect 12466 19472 12478 19506
rect 13254 19472 13266 19506
rect 12466 19460 13266 19472
rect 13947 19506 14747 19518
rect 13947 19472 13959 19506
rect 14735 19472 14747 19506
rect 13947 19460 14747 19472
rect 12466 19248 13266 19260
rect 12466 19214 12478 19248
rect 13254 19214 13266 19248
rect 12466 19202 13266 19214
rect 13947 19248 14747 19260
rect 13947 19214 13959 19248
rect 14735 19214 14747 19248
rect 13947 19202 14747 19214
rect 12466 18990 13266 19002
rect 12466 18956 12478 18990
rect 13254 18956 13266 18990
rect 12466 18944 13266 18956
rect 13947 18990 14747 19002
rect 13947 18956 13959 18990
rect 14735 18956 14747 18990
rect 13947 18944 14747 18956
rect 12466 18732 13266 18744
rect 12466 18698 12478 18732
rect 13254 18698 13266 18732
rect 12466 18686 13266 18698
rect 13947 18732 14747 18744
rect 13947 18698 13959 18732
rect 14735 18698 14747 18732
rect 13947 18686 14747 18698
rect 12466 18474 13266 18486
rect 12466 18440 12478 18474
rect 13254 18440 13266 18474
rect 12466 18428 13266 18440
rect 13947 18474 14747 18486
rect 13947 18440 13959 18474
rect 14735 18440 14747 18474
rect 13947 18428 14747 18440
rect 12466 18216 13266 18228
rect 12466 18182 12478 18216
rect 13254 18182 13266 18216
rect 12466 18170 13266 18182
rect 13947 18216 14747 18228
rect 13947 18182 13959 18216
rect 14735 18182 14747 18216
rect 13947 18170 14747 18182
rect 12466 17958 13266 17970
rect 12466 17924 12478 17958
rect 13254 17924 13266 17958
rect 12466 17912 13266 17924
rect 13947 17958 14747 17970
rect 13947 17924 13959 17958
rect 14735 17924 14747 17958
rect 13947 17912 14747 17924
rect 12466 17700 13266 17712
rect 12466 17666 12478 17700
rect 13254 17666 13266 17700
rect 12466 17654 13266 17666
rect 13947 17700 14747 17712
rect 13947 17666 13959 17700
rect 14735 17666 14747 17700
rect 13947 17654 14747 17666
rect 12466 17442 13266 17454
rect 12466 17408 12478 17442
rect 13254 17408 13266 17442
rect 12466 17396 13266 17408
rect 13947 17442 14747 17454
rect 13947 17408 13959 17442
rect 14735 17408 14747 17442
rect 13947 17396 14747 17408
rect 12466 17184 13266 17196
rect 12466 17150 12478 17184
rect 13254 17150 13266 17184
rect 12466 17138 13266 17150
rect 13947 17184 14747 17196
rect 13947 17150 13959 17184
rect 14735 17150 14747 17184
rect 13947 17138 14747 17150
rect 12466 16926 13266 16938
rect 12466 16892 12478 16926
rect 13254 16892 13266 16926
rect 12466 16880 13266 16892
rect 13947 16926 14747 16938
rect 13947 16892 13959 16926
rect 14735 16892 14747 16926
rect 13947 16880 14747 16892
rect 12466 16668 13266 16680
rect 12466 16634 12478 16668
rect 13254 16634 13266 16668
rect 12466 16622 13266 16634
rect 13947 16668 14747 16680
rect 13947 16634 13959 16668
rect 14735 16634 14747 16668
rect 13947 16622 14747 16634
rect 12466 16410 13266 16422
rect 12466 16376 12478 16410
rect 13254 16376 13266 16410
rect 12466 16364 13266 16376
rect 13947 16410 14747 16422
rect 13947 16376 13959 16410
rect 14735 16376 14747 16410
rect 13947 16364 14747 16376
rect 12466 16152 13266 16164
rect 12466 16118 12478 16152
rect 13254 16118 13266 16152
rect 12466 16106 13266 16118
rect 13947 16152 14747 16164
rect 13947 16118 13959 16152
rect 14735 16118 14747 16152
rect 13947 16106 14747 16118
rect 12466 15894 13266 15906
rect 12466 15860 12478 15894
rect 13254 15860 13266 15894
rect 12466 15848 13266 15860
rect 13947 15894 14747 15906
rect 13947 15860 13959 15894
rect 14735 15860 14747 15894
rect 13947 15848 14747 15860
rect 12466 15636 13266 15648
rect 12466 15602 12478 15636
rect 13254 15602 13266 15636
rect 12466 15590 13266 15602
rect 13947 15636 14747 15648
rect 13947 15602 13959 15636
rect 14735 15602 14747 15636
rect 13947 15590 14747 15602
rect 12466 15378 13266 15390
rect 12466 15344 12478 15378
rect 13254 15344 13266 15378
rect 12466 15332 13266 15344
rect 13947 15378 14747 15390
rect 13947 15344 13959 15378
rect 14735 15344 14747 15378
rect 13947 15332 14747 15344
rect 16084 22375 16284 22387
rect 16084 22341 16096 22375
rect 16272 22341 16284 22375
rect 16084 22329 16284 22341
rect 16084 22117 16284 22129
rect 16084 22083 16096 22117
rect 16272 22083 16284 22117
rect 16084 22071 16284 22083
rect 16084 21859 16284 21871
rect 16084 21825 16096 21859
rect 16272 21825 16284 21859
rect 16084 21813 16284 21825
rect 16084 21601 16284 21613
rect 16084 21567 16096 21601
rect 16272 21567 16284 21601
rect 16084 21555 16284 21567
rect 16084 21343 16284 21355
rect 16084 21309 16096 21343
rect 16272 21309 16284 21343
rect 16084 21297 16284 21309
rect 16084 21085 16284 21097
rect 16084 21051 16096 21085
rect 16272 21051 16284 21085
rect 16084 21039 16284 21051
rect 16084 20827 16284 20839
rect 16084 20793 16096 20827
rect 16272 20793 16284 20827
rect 16084 20781 16284 20793
rect 16084 20569 16284 20581
rect 16084 20535 16096 20569
rect 16272 20535 16284 20569
rect 16084 20523 16284 20535
rect 16084 20311 16284 20323
rect 16084 20277 16096 20311
rect 16272 20277 16284 20311
rect 16084 20265 16284 20277
rect 16084 20053 16284 20065
rect 16084 20019 16096 20053
rect 16272 20019 16284 20053
rect 16084 20007 16284 20019
rect 16084 19795 16284 19807
rect 16084 19761 16096 19795
rect 16272 19761 16284 19795
rect 16084 19749 16284 19761
rect 16084 19537 16284 19549
rect 16084 19503 16096 19537
rect 16272 19503 16284 19537
rect 16084 19491 16284 19503
rect 16084 19279 16284 19291
rect 16084 19245 16096 19279
rect 16272 19245 16284 19279
rect 16084 19233 16284 19245
rect 16084 19021 16284 19033
rect 16084 18987 16096 19021
rect 16272 18987 16284 19021
rect 16084 18975 16284 18987
rect 16084 18763 16284 18775
rect 16084 18729 16096 18763
rect 16272 18729 16284 18763
rect 16084 18717 16284 18729
rect 16084 18505 16284 18517
rect 16084 18471 16096 18505
rect 16272 18471 16284 18505
rect 16084 18459 16284 18471
rect 16084 18247 16284 18259
rect 16084 18213 16096 18247
rect 16272 18213 16284 18247
rect 16084 18201 16284 18213
rect 16084 17989 16284 18001
rect 16084 17955 16096 17989
rect 16272 17955 16284 17989
rect 16084 17943 16284 17955
rect 16084 17731 16284 17743
rect 16084 17697 16096 17731
rect 16272 17697 16284 17731
rect 16084 17685 16284 17697
rect 16084 17473 16284 17485
rect 16084 17439 16096 17473
rect 16272 17439 16284 17473
rect 16084 17427 16284 17439
rect 16084 17215 16284 17227
rect 16084 17181 16096 17215
rect 16272 17181 16284 17215
rect 16084 17169 16284 17181
rect 22654 22750 23754 22762
rect 22654 22716 22666 22750
rect 23742 22716 23754 22750
rect 22654 22704 23754 22716
rect 22654 22392 23754 22404
rect 22654 22358 22666 22392
rect 23742 22358 23754 22392
rect 22654 22346 23754 22358
rect 22654 22034 23754 22046
rect 22654 22000 22666 22034
rect 23742 22000 23754 22034
rect 22654 21988 23754 22000
rect 3101 10185 3901 10197
rect 3101 10151 3113 10185
rect 3889 10151 3901 10185
rect 3101 10139 3901 10151
rect 4582 10185 5382 10197
rect 4582 10151 4594 10185
rect 5370 10151 5382 10185
rect 4582 10139 5382 10151
rect 3101 9927 3901 9939
rect 3101 9893 3113 9927
rect 3889 9893 3901 9927
rect 3101 9881 3901 9893
rect 4582 9927 5382 9939
rect 4582 9893 4594 9927
rect 5370 9893 5382 9927
rect 4582 9881 5382 9893
rect 3101 9669 3901 9681
rect 3101 9635 3113 9669
rect 3889 9635 3901 9669
rect 3101 9623 3901 9635
rect 4582 9669 5382 9681
rect 4582 9635 4594 9669
rect 5370 9635 5382 9669
rect 4582 9623 5382 9635
rect 3101 9411 3901 9423
rect 3101 9377 3113 9411
rect 3889 9377 3901 9411
rect 3101 9365 3901 9377
rect 4582 9411 5382 9423
rect 4582 9377 4594 9411
rect 5370 9377 5382 9411
rect 4582 9365 5382 9377
rect 3101 9153 3901 9165
rect 3101 9119 3113 9153
rect 3889 9119 3901 9153
rect 3101 9107 3901 9119
rect 4582 9153 5382 9165
rect 4582 9119 4594 9153
rect 5370 9119 5382 9153
rect 4582 9107 5382 9119
rect 3101 8895 3901 8907
rect 3101 8861 3113 8895
rect 3889 8861 3901 8895
rect 3101 8849 3901 8861
rect 4582 8895 5382 8907
rect 4582 8861 4594 8895
rect 5370 8861 5382 8895
rect 4582 8849 5382 8861
rect 3101 8637 3901 8649
rect 3101 8603 3113 8637
rect 3889 8603 3901 8637
rect 3101 8591 3901 8603
rect 4582 8637 5382 8649
rect 4582 8603 4594 8637
rect 5370 8603 5382 8637
rect 4582 8591 5382 8603
rect 3101 8379 3901 8391
rect 3101 8345 3113 8379
rect 3889 8345 3901 8379
rect 3101 8333 3901 8345
rect 4582 8379 5382 8391
rect 4582 8345 4594 8379
rect 5370 8345 5382 8379
rect 4582 8333 5382 8345
rect 3101 8121 3901 8133
rect 3101 8087 3113 8121
rect 3889 8087 3901 8121
rect 3101 8075 3901 8087
rect 4582 8121 5382 8133
rect 4582 8087 4594 8121
rect 5370 8087 5382 8121
rect 4582 8075 5382 8087
rect 3101 7863 3901 7875
rect 3101 7829 3113 7863
rect 3889 7829 3901 7863
rect 3101 7817 3901 7829
rect 4582 7863 5382 7875
rect 4582 7829 4594 7863
rect 5370 7829 5382 7863
rect 4582 7817 5382 7829
rect 3101 7605 3901 7617
rect 3101 7571 3113 7605
rect 3889 7571 3901 7605
rect 3101 7559 3901 7571
rect 4582 7605 5382 7617
rect 4582 7571 4594 7605
rect 5370 7571 5382 7605
rect 4582 7559 5382 7571
rect 3101 7347 3901 7359
rect 3101 7313 3113 7347
rect 3889 7313 3901 7347
rect 3101 7301 3901 7313
rect 4582 7347 5382 7359
rect 4582 7313 4594 7347
rect 5370 7313 5382 7347
rect 4582 7301 5382 7313
rect 3101 7089 3901 7101
rect 3101 7055 3113 7089
rect 3889 7055 3901 7089
rect 3101 7043 3901 7055
rect 4582 7089 5382 7101
rect 4582 7055 4594 7089
rect 5370 7055 5382 7089
rect 4582 7043 5382 7055
rect 3101 6831 3901 6843
rect 3101 6797 3113 6831
rect 3889 6797 3901 6831
rect 3101 6785 3901 6797
rect 4582 6831 5382 6843
rect 4582 6797 4594 6831
rect 5370 6797 5382 6831
rect 4582 6785 5382 6797
rect 3101 6573 3901 6585
rect 3101 6539 3113 6573
rect 3889 6539 3901 6573
rect 3101 6527 3901 6539
rect 4582 6573 5382 6585
rect 4582 6539 4594 6573
rect 5370 6539 5382 6573
rect 4582 6527 5382 6539
rect 3101 6315 3901 6327
rect 3101 6281 3113 6315
rect 3889 6281 3901 6315
rect 3101 6269 3901 6281
rect 4582 6315 5382 6327
rect 4582 6281 4594 6315
rect 5370 6281 5382 6315
rect 4582 6269 5382 6281
rect 3101 6057 3901 6069
rect 3101 6023 3113 6057
rect 3889 6023 3901 6057
rect 3101 6011 3901 6023
rect 4582 6057 5382 6069
rect 4582 6023 4594 6057
rect 5370 6023 5382 6057
rect 4582 6011 5382 6023
rect 3101 5799 3901 5811
rect 3101 5765 3113 5799
rect 3889 5765 3901 5799
rect 3101 5753 3901 5765
rect 4582 5799 5382 5811
rect 4582 5765 4594 5799
rect 5370 5765 5382 5799
rect 4582 5753 5382 5765
rect 3101 5541 3901 5553
rect 3101 5507 3113 5541
rect 3889 5507 3901 5541
rect 3101 5495 3901 5507
rect 4582 5541 5382 5553
rect 4582 5507 4594 5541
rect 5370 5507 5382 5541
rect 4582 5495 5382 5507
rect 3101 5283 3901 5295
rect 3101 5249 3113 5283
rect 3889 5249 3901 5283
rect 3101 5237 3901 5249
rect 4582 5283 5382 5295
rect 4582 5249 4594 5283
rect 5370 5249 5382 5283
rect 4582 5237 5382 5249
rect 3101 5025 3901 5037
rect 3101 4991 3113 5025
rect 3889 4991 3901 5025
rect 3101 4979 3901 4991
rect 4582 5025 5382 5037
rect 4582 4991 4594 5025
rect 5370 4991 5382 5025
rect 4582 4979 5382 4991
rect 3101 4767 3901 4779
rect 3101 4733 3113 4767
rect 3889 4733 3901 4767
rect 3101 4721 3901 4733
rect 4582 4767 5382 4779
rect 4582 4733 4594 4767
rect 5370 4733 5382 4767
rect 4582 4721 5382 4733
rect 3101 4509 3901 4521
rect 3101 4475 3113 4509
rect 3889 4475 3901 4509
rect 3101 4463 3901 4475
rect 4582 4509 5382 4521
rect 4582 4475 4594 4509
rect 5370 4475 5382 4509
rect 4582 4463 5382 4475
rect 3101 4251 3901 4263
rect 3101 4217 3113 4251
rect 3889 4217 3901 4251
rect 3101 4205 3901 4217
rect 4582 4251 5382 4263
rect 4582 4217 4594 4251
rect 5370 4217 5382 4251
rect 4582 4205 5382 4217
rect 3101 3993 3901 4005
rect 3101 3959 3113 3993
rect 3889 3959 3901 3993
rect 3101 3947 3901 3959
rect 4582 3993 5382 4005
rect 4582 3959 4594 3993
rect 5370 3959 5382 3993
rect 4582 3947 5382 3959
rect 6719 8249 6919 8261
rect 6719 8215 6731 8249
rect 6907 8215 6919 8249
rect 6719 8203 6919 8215
rect 6719 7991 6919 8003
rect 6719 7957 6731 7991
rect 6907 7957 6919 7991
rect 6719 7945 6919 7957
rect 6719 7733 6919 7745
rect 6719 7699 6731 7733
rect 6907 7699 6919 7733
rect 6719 7687 6919 7699
rect 6719 7475 6919 7487
rect 6719 7441 6731 7475
rect 6907 7441 6919 7475
rect 6719 7429 6919 7441
rect 6719 7217 6919 7229
rect 6719 7183 6731 7217
rect 6907 7183 6919 7217
rect 6719 7171 6919 7183
rect 6719 6959 6919 6971
rect 6719 6925 6731 6959
rect 6907 6925 6919 6959
rect 6719 6913 6919 6925
rect 6719 6701 6919 6713
rect 6719 6667 6731 6701
rect 6907 6667 6919 6701
rect 6719 6655 6919 6667
rect 6719 6443 6919 6455
rect 6719 6409 6731 6443
rect 6907 6409 6919 6443
rect 6719 6397 6919 6409
rect 6719 6185 6919 6197
rect 6719 6151 6731 6185
rect 6907 6151 6919 6185
rect 6719 6139 6919 6151
rect 6719 5927 6919 5939
rect 6719 5893 6731 5927
rect 6907 5893 6919 5927
rect 6719 5881 6919 5893
rect 6719 5669 6919 5681
rect 6719 5635 6731 5669
rect 6907 5635 6919 5669
rect 6719 5623 6919 5635
rect 6719 5411 6919 5423
rect 6719 5377 6731 5411
rect 6907 5377 6919 5411
rect 6719 5365 6919 5377
rect 6719 5153 6919 5165
rect 6719 5119 6731 5153
rect 6907 5119 6919 5153
rect 6719 5107 6919 5119
rect 6719 4895 6919 4907
rect 6719 4861 6731 4895
rect 6907 4861 6919 4895
rect 6719 4849 6919 4861
rect 6719 4637 6919 4649
rect 6719 4603 6731 4637
rect 6907 4603 6919 4637
rect 6719 4591 6919 4603
rect 6719 4379 6919 4391
rect 6719 4345 6731 4379
rect 6907 4345 6919 4379
rect 6719 4333 6919 4345
rect 6719 4121 6919 4133
rect 6719 4087 6731 4121
rect 6907 4087 6919 4121
rect 6719 4075 6919 4087
rect 6719 3863 6919 3875
rect 6719 3829 6731 3863
rect 6907 3829 6919 3863
rect 6719 3817 6919 3829
rect 6719 3605 6919 3617
rect 6719 3571 6731 3605
rect 6907 3571 6919 3605
rect 6719 3559 6919 3571
rect 6719 3347 6919 3359
rect 6719 3313 6731 3347
rect 6907 3313 6919 3347
rect 6719 3301 6919 3313
rect 6719 3089 6919 3101
rect 6719 3055 6731 3089
rect 6907 3055 6919 3089
rect 6719 3043 6919 3055
rect 18046 7269 18646 7281
rect 18046 7235 18058 7269
rect 18634 7235 18646 7269
rect 18046 7223 18646 7235
rect 18046 6211 18646 6223
rect 18046 6177 18058 6211
rect 18634 6177 18646 6211
rect 18046 6165 18646 6177
rect 19373 8782 19431 8794
rect 19373 7606 19385 8782
rect 19419 7606 19431 8782
rect 19373 7594 19431 7606
rect 21831 8782 21889 8794
rect 21831 7606 21843 8782
rect 21877 7606 21889 8782
rect 21831 7594 21889 7606
rect 24289 8782 24347 8794
rect 24289 7606 24301 8782
rect 24335 7606 24347 8782
rect 24289 7594 24347 7606
rect 19372 6907 19430 6919
rect 19372 5731 19384 6907
rect 19418 5731 19430 6907
rect 19372 5719 19430 5731
rect 21830 6907 21888 6919
rect 21830 5731 21842 6907
rect 21876 5731 21888 6907
rect 21830 5719 21888 5731
rect 24288 6907 24346 6919
rect 24288 5731 24300 6907
rect 24334 5731 24346 6907
rect 24288 5719 24346 5731
<< pdiff >>
rect 3654 30440 3712 30452
rect 3654 30104 3666 30440
rect 3700 30104 3712 30440
rect 3654 30092 3712 30104
rect 7312 30440 7370 30452
rect 7312 30104 7324 30440
rect 7358 30104 7370 30440
rect 7312 30092 7370 30104
rect 10970 30440 11028 30452
rect 10970 30104 10982 30440
rect 11016 30104 11028 30440
rect 10970 30092 11028 30104
rect 3654 29952 3712 29964
rect 3654 29616 3666 29952
rect 3700 29616 3712 29952
rect 3654 29604 3712 29616
rect 7312 29952 7370 29964
rect 7312 29616 7324 29952
rect 7358 29616 7370 29952
rect 7312 29604 7370 29616
rect 10970 29952 11028 29964
rect 10970 29616 10982 29952
rect 11016 29616 11028 29952
rect 10970 29604 11028 29616
rect 12126 32516 12184 32528
rect 12126 29540 12138 32516
rect 12172 29540 12184 32516
rect 12126 29528 12184 29540
rect 12564 32516 12622 32528
rect 12564 29540 12576 32516
rect 12610 29540 12622 32516
rect 12564 29528 12622 29540
rect 13002 32516 13060 32528
rect 13002 29540 13014 32516
rect 13048 29540 13060 32516
rect 13002 29528 13060 29540
rect 13440 32516 13498 32528
rect 13440 29540 13452 32516
rect 13486 29540 13498 32516
rect 13440 29528 13498 29540
rect 13878 32516 13936 32528
rect 13878 29540 13890 32516
rect 13924 29540 13936 32516
rect 13878 29528 13936 29540
rect 12126 28539 12184 28551
rect 12126 25563 12138 28539
rect 12172 25563 12184 28539
rect 12126 25551 12184 25563
rect 12564 28539 12622 28551
rect 12564 25563 12576 28539
rect 12610 25563 12622 28539
rect 12564 25551 12622 25563
rect 13002 28539 13060 28551
rect 13002 25563 13014 28539
rect 13048 25563 13060 28539
rect 13002 25551 13060 25563
rect 13440 28539 13498 28551
rect 13440 25563 13452 28539
rect 13486 25563 13498 28539
rect 13440 25551 13498 25563
rect 13878 28539 13936 28551
rect 13878 25563 13890 28539
rect 13924 25563 13936 28539
rect 13878 25551 13936 25563
rect 16955 26985 17013 26997
rect 16955 25609 16967 26985
rect 17001 25609 17013 26985
rect 16955 25597 17013 25609
rect 17373 26985 17431 26997
rect 17373 25609 17385 26985
rect 17419 25609 17431 26985
rect 17373 25597 17431 25609
rect 17791 26985 17849 26997
rect 17791 25609 17803 26985
rect 17837 25609 17849 26985
rect 17791 25597 17849 25609
rect 18209 26985 18267 26997
rect 18209 25609 18221 26985
rect 18255 25609 18267 26985
rect 18209 25597 18267 25609
rect 18627 26985 18685 26997
rect 18627 25609 18639 26985
rect 18673 25609 18685 26985
rect 18627 25597 18685 25609
rect 21048 27530 21106 27542
rect 21048 27054 21060 27530
rect 21094 27054 21106 27530
rect 21048 27042 21106 27054
rect 22106 27530 22164 27542
rect 22106 27054 22118 27530
rect 22152 27054 22164 27530
rect 22106 27042 22164 27054
rect 23164 27530 23222 27542
rect 23164 27054 23176 27530
rect 23210 27054 23222 27530
rect 23164 27042 23222 27054
rect 24222 27530 24280 27542
rect 24222 27054 24234 27530
rect 24268 27054 24280 27530
rect 24222 27042 24280 27054
rect 25280 27530 25338 27542
rect 25280 27054 25292 27530
rect 25326 27054 25338 27530
rect 25280 27042 25338 27054
rect 21048 26368 21106 26380
rect 21048 25892 21060 26368
rect 21094 25892 21106 26368
rect 21048 25880 21106 25892
rect 22106 26368 22164 26380
rect 22106 25892 22118 26368
rect 22152 25892 22164 26368
rect 22106 25880 22164 25892
rect 23164 26368 23222 26380
rect 23164 25892 23176 26368
rect 23210 25892 23222 26368
rect 23164 25880 23222 25892
rect 24222 26368 24280 26380
rect 24222 25892 24234 26368
rect 24268 25892 24280 26368
rect 24222 25880 24280 25892
rect 25280 26368 25338 26380
rect 25280 25892 25292 26368
rect 25326 25892 25338 26368
rect 25280 25880 25338 25892
rect 25381 24965 25439 24977
rect 25381 24469 25393 24965
rect 25427 24469 25439 24965
rect 25381 24457 25439 24469
rect 25509 24965 25567 24977
rect 25509 24469 25521 24965
rect 25555 24469 25567 24965
rect 25509 24457 25567 24469
rect 25737 24965 25795 24977
rect 25737 24469 25749 24965
rect 25783 24469 25795 24965
rect 25737 24457 25795 24469
rect 25865 24965 25923 24977
rect 25865 24469 25877 24965
rect 25911 24469 25923 24965
rect 25865 24457 25923 24469
rect 16871 22440 17071 22452
rect 16871 22406 16883 22440
rect 17059 22406 17071 22440
rect 16871 22394 17071 22406
rect 16871 21982 17071 21994
rect 16871 21948 16883 21982
rect 17059 21948 17071 21982
rect 16871 21936 17071 21948
rect 16871 21859 17071 21871
rect 16871 21825 16883 21859
rect 17059 21825 17071 21859
rect 16871 21813 17071 21825
rect 16871 21401 17071 21413
rect 16871 21367 16883 21401
rect 17059 21367 17071 21401
rect 16871 21355 17071 21367
rect 16871 20569 17071 20581
rect 16871 20535 16883 20569
rect 17059 20535 17071 20569
rect 16871 20523 17071 20535
rect 16871 20111 17071 20123
rect 16871 20077 16883 20111
rect 17059 20077 17071 20111
rect 16871 20065 17071 20077
rect 16871 19279 17071 19291
rect 16871 19245 16883 19279
rect 17059 19245 17071 19279
rect 16871 19233 17071 19245
rect 16871 18821 17071 18833
rect 16871 18787 16883 18821
rect 17059 18787 17071 18821
rect 16871 18775 17071 18787
rect 16871 17989 17071 18001
rect 16871 17955 16883 17989
rect 17059 17955 17071 17989
rect 16871 17943 17071 17955
rect 16871 17531 17071 17543
rect 16871 17497 16883 17531
rect 17059 17497 17071 17531
rect 16871 17485 17071 17497
rect 16871 16901 17071 16913
rect 16871 16867 16883 16901
rect 17059 16867 17071 16901
rect 16871 16855 17071 16867
rect 15540 16036 16220 16088
rect 15540 16002 15592 16036
rect 15626 16002 15682 16036
rect 15716 16002 15772 16036
rect 15806 16002 15862 16036
rect 15896 16002 15952 16036
rect 15986 16002 16042 16036
rect 16076 16002 16132 16036
rect 16166 16002 16220 16036
rect 15540 15946 16220 16002
rect 15540 15912 15592 15946
rect 15626 15912 15682 15946
rect 15716 15912 15772 15946
rect 15806 15912 15862 15946
rect 15896 15912 15952 15946
rect 15986 15912 16042 15946
rect 16076 15912 16132 15946
rect 16166 15912 16220 15946
rect 15540 15856 16220 15912
rect 15540 15822 15592 15856
rect 15626 15822 15682 15856
rect 15716 15822 15772 15856
rect 15806 15822 15862 15856
rect 15896 15822 15952 15856
rect 15986 15822 16042 15856
rect 16076 15822 16132 15856
rect 16166 15822 16220 15856
rect 15540 15766 16220 15822
rect 15540 15732 15592 15766
rect 15626 15732 15682 15766
rect 15716 15732 15772 15766
rect 15806 15732 15862 15766
rect 15896 15732 15952 15766
rect 15986 15732 16042 15766
rect 16076 15732 16132 15766
rect 16166 15732 16220 15766
rect 15540 15676 16220 15732
rect 15540 15642 15592 15676
rect 15626 15642 15682 15676
rect 15716 15642 15772 15676
rect 15806 15642 15862 15676
rect 15896 15642 15952 15676
rect 15986 15642 16042 15676
rect 16076 15642 16132 15676
rect 16166 15642 16220 15676
rect 15540 15586 16220 15642
rect 15540 15552 15592 15586
rect 15626 15552 15682 15586
rect 15716 15552 15772 15586
rect 15806 15552 15862 15586
rect 15896 15552 15952 15586
rect 15986 15552 16042 15586
rect 16076 15552 16132 15586
rect 16166 15552 16220 15586
rect 15540 15496 16220 15552
rect 15540 15462 15592 15496
rect 15626 15462 15682 15496
rect 15716 15462 15772 15496
rect 15806 15462 15862 15496
rect 15896 15462 15952 15496
rect 15986 15462 16042 15496
rect 16076 15462 16132 15496
rect 16166 15462 16220 15496
rect 15540 15408 16220 15462
rect 16871 16643 17071 16655
rect 16871 16609 16883 16643
rect 17059 16609 17071 16643
rect 16871 16597 17071 16609
rect 16871 16385 17071 16397
rect 16871 16351 16883 16385
rect 17059 16351 17071 16385
rect 16871 16339 17071 16351
rect 16871 16176 16971 16188
rect 16871 16142 16883 16176
rect 16959 16142 16971 16176
rect 16871 16130 16971 16142
rect 16871 15718 16971 15730
rect 16871 15684 16883 15718
rect 16959 15684 16971 15718
rect 16871 15672 16971 15684
rect 16871 15260 16971 15272
rect 16871 15226 16883 15260
rect 16959 15226 16971 15260
rect 16871 15214 16971 15226
rect 6175 10067 6855 10121
rect 6175 10033 6227 10067
rect 6261 10033 6317 10067
rect 6351 10033 6407 10067
rect 6441 10033 6497 10067
rect 6531 10033 6587 10067
rect 6621 10033 6677 10067
rect 6711 10033 6767 10067
rect 6801 10033 6855 10067
rect 6175 9977 6855 10033
rect 6175 9943 6227 9977
rect 6261 9943 6317 9977
rect 6351 9943 6407 9977
rect 6441 9943 6497 9977
rect 6531 9943 6587 9977
rect 6621 9943 6677 9977
rect 6711 9943 6767 9977
rect 6801 9943 6855 9977
rect 6175 9887 6855 9943
rect 6175 9853 6227 9887
rect 6261 9853 6317 9887
rect 6351 9853 6407 9887
rect 6441 9853 6497 9887
rect 6531 9853 6587 9887
rect 6621 9853 6677 9887
rect 6711 9853 6767 9887
rect 6801 9853 6855 9887
rect 6175 9797 6855 9853
rect 6175 9763 6227 9797
rect 6261 9763 6317 9797
rect 6351 9763 6407 9797
rect 6441 9763 6497 9797
rect 6531 9763 6587 9797
rect 6621 9763 6677 9797
rect 6711 9763 6767 9797
rect 6801 9763 6855 9797
rect 6175 9707 6855 9763
rect 6175 9673 6227 9707
rect 6261 9673 6317 9707
rect 6351 9673 6407 9707
rect 6441 9673 6497 9707
rect 6531 9673 6587 9707
rect 6621 9673 6677 9707
rect 6711 9673 6767 9707
rect 6801 9673 6855 9707
rect 6175 9617 6855 9673
rect 6175 9583 6227 9617
rect 6261 9583 6317 9617
rect 6351 9583 6407 9617
rect 6441 9583 6497 9617
rect 6531 9583 6587 9617
rect 6621 9583 6677 9617
rect 6711 9583 6767 9617
rect 6801 9583 6855 9617
rect 6175 9527 6855 9583
rect 6175 9493 6227 9527
rect 6261 9493 6317 9527
rect 6351 9493 6407 9527
rect 6441 9493 6497 9527
rect 6531 9493 6587 9527
rect 6621 9493 6677 9527
rect 6711 9493 6767 9527
rect 6801 9493 6855 9527
rect 6175 9441 6855 9493
rect 7506 10303 7606 10315
rect 7506 10269 7518 10303
rect 7594 10269 7606 10303
rect 7506 10257 7606 10269
rect 7506 9845 7606 9857
rect 7506 9811 7518 9845
rect 7594 9811 7606 9845
rect 7506 9799 7606 9811
rect 7506 9387 7606 9399
rect 7506 9353 7518 9387
rect 7594 9353 7606 9387
rect 7506 9341 7606 9353
rect 7506 9178 7706 9190
rect 7506 9144 7518 9178
rect 7694 9144 7706 9178
rect 7506 9132 7706 9144
rect 7506 8920 7706 8932
rect 7506 8886 7518 8920
rect 7694 8886 7706 8920
rect 7506 8874 7706 8886
rect 7506 8662 7706 8674
rect 7506 8628 7518 8662
rect 7694 8628 7706 8662
rect 7506 8616 7706 8628
rect 18163 10654 18221 10666
rect 18163 10318 18175 10654
rect 18209 10318 18221 10654
rect 18163 10306 18221 10318
rect 21821 10654 21879 10666
rect 21821 10318 21833 10654
rect 21867 10318 21879 10654
rect 21821 10306 21879 10318
rect 25479 10654 25537 10666
rect 25479 10318 25491 10654
rect 25525 10318 25537 10654
rect 25479 10306 25537 10318
rect 18163 10166 18221 10178
rect 18163 9830 18175 10166
rect 18209 9830 18221 10166
rect 18163 9818 18221 9830
rect 21821 10166 21879 10178
rect 21821 9830 21833 10166
rect 21867 9830 21879 10166
rect 21821 9818 21879 9830
rect 25479 10166 25537 10178
rect 25479 9830 25491 10166
rect 25525 9830 25537 10166
rect 25479 9818 25537 9830
rect 7506 7933 7706 7945
rect 7506 7899 7518 7933
rect 7694 7899 7706 7933
rect 7506 7887 7706 7899
rect 7506 7475 7706 7487
rect 7506 7441 7518 7475
rect 7694 7441 7706 7475
rect 7506 7429 7706 7441
rect 7506 6643 7706 6655
rect 7506 6609 7518 6643
rect 7694 6609 7706 6643
rect 7506 6597 7706 6609
rect 7506 6185 7706 6197
rect 7506 6151 7518 6185
rect 7694 6151 7706 6185
rect 7506 6139 7706 6151
rect 7506 5353 7706 5365
rect 7506 5319 7518 5353
rect 7694 5319 7706 5353
rect 7506 5307 7706 5319
rect 7506 4895 7706 4907
rect 7506 4861 7518 4895
rect 7694 4861 7706 4895
rect 7506 4849 7706 4861
rect 7506 4063 7706 4075
rect 7506 4029 7518 4063
rect 7694 4029 7706 4063
rect 7506 4017 7706 4029
rect 7506 3605 7706 3617
rect 7506 3571 7518 3605
rect 7694 3571 7706 3605
rect 7506 3559 7706 3571
rect 7506 3482 7706 3494
rect 7506 3448 7518 3482
rect 7694 3448 7706 3482
rect 7506 3436 7706 3448
rect 7506 3024 7706 3036
rect 7506 2990 7518 3024
rect 7694 2990 7706 3024
rect 7506 2978 7706 2990
<< ndiffc >>
rect 3549 27021 4125 27055
rect 3549 25963 4125 25997
rect 4876 27392 4910 28568
rect 7334 27392 7368 28568
rect 9792 27392 9826 28568
rect 4875 25517 4909 26693
rect 7333 25517 7367 26693
rect 9791 25517 9825 26693
rect 12148 24237 12182 24513
rect 14086 24237 14120 24513
rect 16024 24237 16058 24513
rect 17962 24237 17996 24513
rect 19900 24237 19934 24513
rect 12148 23827 12182 24103
rect 14086 23827 14120 24103
rect 16024 23827 16058 24103
rect 17962 23827 17996 24103
rect 19900 23827 19934 24103
rect 22245 24507 22279 25083
rect 22703 24507 22737 25083
rect 23161 24507 23195 25083
rect 23619 24507 23653 25083
rect 24077 24507 24111 25083
rect 22245 23300 22279 23876
rect 22703 23300 22737 23876
rect 23161 23300 23195 23876
rect 23619 23300 23653 23876
rect 24077 23300 24111 23876
rect 25433 23784 25467 23960
rect 25521 23784 25555 23960
rect 25789 23784 25823 23960
rect 25877 23784 25911 23960
rect 12478 21536 13254 21570
rect 13959 21536 14735 21570
rect 12478 21278 13254 21312
rect 13959 21278 14735 21312
rect 12478 21020 13254 21054
rect 13959 21020 14735 21054
rect 12478 20762 13254 20796
rect 13959 20762 14735 20796
rect 12478 20504 13254 20538
rect 13959 20504 14735 20538
rect 12478 20246 13254 20280
rect 13959 20246 14735 20280
rect 12478 19988 13254 20022
rect 13959 19988 14735 20022
rect 12478 19730 13254 19764
rect 13959 19730 14735 19764
rect 12478 19472 13254 19506
rect 13959 19472 14735 19506
rect 12478 19214 13254 19248
rect 13959 19214 14735 19248
rect 12478 18956 13254 18990
rect 13959 18956 14735 18990
rect 12478 18698 13254 18732
rect 13959 18698 14735 18732
rect 12478 18440 13254 18474
rect 13959 18440 14735 18474
rect 12478 18182 13254 18216
rect 13959 18182 14735 18216
rect 12478 17924 13254 17958
rect 13959 17924 14735 17958
rect 12478 17666 13254 17700
rect 13959 17666 14735 17700
rect 12478 17408 13254 17442
rect 13959 17408 14735 17442
rect 12478 17150 13254 17184
rect 13959 17150 14735 17184
rect 12478 16892 13254 16926
rect 13959 16892 14735 16926
rect 12478 16634 13254 16668
rect 13959 16634 14735 16668
rect 12478 16376 13254 16410
rect 13959 16376 14735 16410
rect 12478 16118 13254 16152
rect 13959 16118 14735 16152
rect 12478 15860 13254 15894
rect 13959 15860 14735 15894
rect 12478 15602 13254 15636
rect 13959 15602 14735 15636
rect 12478 15344 13254 15378
rect 13959 15344 14735 15378
rect 16096 22341 16272 22375
rect 16096 22083 16272 22117
rect 16096 21825 16272 21859
rect 16096 21567 16272 21601
rect 16096 21309 16272 21343
rect 16096 21051 16272 21085
rect 16096 20793 16272 20827
rect 16096 20535 16272 20569
rect 16096 20277 16272 20311
rect 16096 20019 16272 20053
rect 16096 19761 16272 19795
rect 16096 19503 16272 19537
rect 16096 19245 16272 19279
rect 16096 18987 16272 19021
rect 16096 18729 16272 18763
rect 16096 18471 16272 18505
rect 16096 18213 16272 18247
rect 16096 17955 16272 17989
rect 16096 17697 16272 17731
rect 16096 17439 16272 17473
rect 16096 17181 16272 17215
rect 22666 22716 23742 22750
rect 22666 22358 23742 22392
rect 22666 22000 23742 22034
rect 3113 10151 3889 10185
rect 4594 10151 5370 10185
rect 3113 9893 3889 9927
rect 4594 9893 5370 9927
rect 3113 9635 3889 9669
rect 4594 9635 5370 9669
rect 3113 9377 3889 9411
rect 4594 9377 5370 9411
rect 3113 9119 3889 9153
rect 4594 9119 5370 9153
rect 3113 8861 3889 8895
rect 4594 8861 5370 8895
rect 3113 8603 3889 8637
rect 4594 8603 5370 8637
rect 3113 8345 3889 8379
rect 4594 8345 5370 8379
rect 3113 8087 3889 8121
rect 4594 8087 5370 8121
rect 3113 7829 3889 7863
rect 4594 7829 5370 7863
rect 3113 7571 3889 7605
rect 4594 7571 5370 7605
rect 3113 7313 3889 7347
rect 4594 7313 5370 7347
rect 3113 7055 3889 7089
rect 4594 7055 5370 7089
rect 3113 6797 3889 6831
rect 4594 6797 5370 6831
rect 3113 6539 3889 6573
rect 4594 6539 5370 6573
rect 3113 6281 3889 6315
rect 4594 6281 5370 6315
rect 3113 6023 3889 6057
rect 4594 6023 5370 6057
rect 3113 5765 3889 5799
rect 4594 5765 5370 5799
rect 3113 5507 3889 5541
rect 4594 5507 5370 5541
rect 3113 5249 3889 5283
rect 4594 5249 5370 5283
rect 3113 4991 3889 5025
rect 4594 4991 5370 5025
rect 3113 4733 3889 4767
rect 4594 4733 5370 4767
rect 3113 4475 3889 4509
rect 4594 4475 5370 4509
rect 3113 4217 3889 4251
rect 4594 4217 5370 4251
rect 3113 3959 3889 3993
rect 4594 3959 5370 3993
rect 6731 8215 6907 8249
rect 6731 7957 6907 7991
rect 6731 7699 6907 7733
rect 6731 7441 6907 7475
rect 6731 7183 6907 7217
rect 6731 6925 6907 6959
rect 6731 6667 6907 6701
rect 6731 6409 6907 6443
rect 6731 6151 6907 6185
rect 6731 5893 6907 5927
rect 6731 5635 6907 5669
rect 6731 5377 6907 5411
rect 6731 5119 6907 5153
rect 6731 4861 6907 4895
rect 6731 4603 6907 4637
rect 6731 4345 6907 4379
rect 6731 4087 6907 4121
rect 6731 3829 6907 3863
rect 6731 3571 6907 3605
rect 6731 3313 6907 3347
rect 6731 3055 6907 3089
rect 18058 7235 18634 7269
rect 18058 6177 18634 6211
rect 19385 7606 19419 8782
rect 21843 7606 21877 8782
rect 24301 7606 24335 8782
rect 19384 5731 19418 6907
rect 21842 5731 21876 6907
rect 24300 5731 24334 6907
<< pdiffc >>
rect 3666 30104 3700 30440
rect 7324 30104 7358 30440
rect 10982 30104 11016 30440
rect 3666 29616 3700 29952
rect 7324 29616 7358 29952
rect 10982 29616 11016 29952
rect 12138 29540 12172 32516
rect 12576 29540 12610 32516
rect 13014 29540 13048 32516
rect 13452 29540 13486 32516
rect 13890 29540 13924 32516
rect 12138 25563 12172 28539
rect 12576 25563 12610 28539
rect 13014 25563 13048 28539
rect 13452 25563 13486 28539
rect 13890 25563 13924 28539
rect 16967 25609 17001 26985
rect 17385 25609 17419 26985
rect 17803 25609 17837 26985
rect 18221 25609 18255 26985
rect 18639 25609 18673 26985
rect 21060 27054 21094 27530
rect 22118 27054 22152 27530
rect 23176 27054 23210 27530
rect 24234 27054 24268 27530
rect 25292 27054 25326 27530
rect 21060 25892 21094 26368
rect 22118 25892 22152 26368
rect 23176 25892 23210 26368
rect 24234 25892 24268 26368
rect 25292 25892 25326 26368
rect 25393 24469 25427 24965
rect 25521 24469 25555 24965
rect 25749 24469 25783 24965
rect 25877 24469 25911 24965
rect 16883 22406 17059 22440
rect 16883 21948 17059 21982
rect 16883 21825 17059 21859
rect 16883 21367 17059 21401
rect 16883 20535 17059 20569
rect 16883 20077 17059 20111
rect 16883 19245 17059 19279
rect 16883 18787 17059 18821
rect 16883 17955 17059 17989
rect 16883 17497 17059 17531
rect 16883 16867 17059 16901
rect 15592 16002 15626 16036
rect 15682 16002 15716 16036
rect 15772 16002 15806 16036
rect 15862 16002 15896 16036
rect 15952 16002 15986 16036
rect 16042 16002 16076 16036
rect 16132 16002 16166 16036
rect 15592 15912 15626 15946
rect 15682 15912 15716 15946
rect 15772 15912 15806 15946
rect 15862 15912 15896 15946
rect 15952 15912 15986 15946
rect 16042 15912 16076 15946
rect 16132 15912 16166 15946
rect 15592 15822 15626 15856
rect 15682 15822 15716 15856
rect 15772 15822 15806 15856
rect 15862 15822 15896 15856
rect 15952 15822 15986 15856
rect 16042 15822 16076 15856
rect 16132 15822 16166 15856
rect 15592 15732 15626 15766
rect 15682 15732 15716 15766
rect 15772 15732 15806 15766
rect 15862 15732 15896 15766
rect 15952 15732 15986 15766
rect 16042 15732 16076 15766
rect 16132 15732 16166 15766
rect 15592 15642 15626 15676
rect 15682 15642 15716 15676
rect 15772 15642 15806 15676
rect 15862 15642 15896 15676
rect 15952 15642 15986 15676
rect 16042 15642 16076 15676
rect 16132 15642 16166 15676
rect 15592 15552 15626 15586
rect 15682 15552 15716 15586
rect 15772 15552 15806 15586
rect 15862 15552 15896 15586
rect 15952 15552 15986 15586
rect 16042 15552 16076 15586
rect 16132 15552 16166 15586
rect 15592 15462 15626 15496
rect 15682 15462 15716 15496
rect 15772 15462 15806 15496
rect 15862 15462 15896 15496
rect 15952 15462 15986 15496
rect 16042 15462 16076 15496
rect 16132 15462 16166 15496
rect 16883 16609 17059 16643
rect 16883 16351 17059 16385
rect 16883 16142 16959 16176
rect 16883 15684 16959 15718
rect 16883 15226 16959 15260
rect 6227 10033 6261 10067
rect 6317 10033 6351 10067
rect 6407 10033 6441 10067
rect 6497 10033 6531 10067
rect 6587 10033 6621 10067
rect 6677 10033 6711 10067
rect 6767 10033 6801 10067
rect 6227 9943 6261 9977
rect 6317 9943 6351 9977
rect 6407 9943 6441 9977
rect 6497 9943 6531 9977
rect 6587 9943 6621 9977
rect 6677 9943 6711 9977
rect 6767 9943 6801 9977
rect 6227 9853 6261 9887
rect 6317 9853 6351 9887
rect 6407 9853 6441 9887
rect 6497 9853 6531 9887
rect 6587 9853 6621 9887
rect 6677 9853 6711 9887
rect 6767 9853 6801 9887
rect 6227 9763 6261 9797
rect 6317 9763 6351 9797
rect 6407 9763 6441 9797
rect 6497 9763 6531 9797
rect 6587 9763 6621 9797
rect 6677 9763 6711 9797
rect 6767 9763 6801 9797
rect 6227 9673 6261 9707
rect 6317 9673 6351 9707
rect 6407 9673 6441 9707
rect 6497 9673 6531 9707
rect 6587 9673 6621 9707
rect 6677 9673 6711 9707
rect 6767 9673 6801 9707
rect 6227 9583 6261 9617
rect 6317 9583 6351 9617
rect 6407 9583 6441 9617
rect 6497 9583 6531 9617
rect 6587 9583 6621 9617
rect 6677 9583 6711 9617
rect 6767 9583 6801 9617
rect 6227 9493 6261 9527
rect 6317 9493 6351 9527
rect 6407 9493 6441 9527
rect 6497 9493 6531 9527
rect 6587 9493 6621 9527
rect 6677 9493 6711 9527
rect 6767 9493 6801 9527
rect 7518 10269 7594 10303
rect 7518 9811 7594 9845
rect 7518 9353 7594 9387
rect 7518 9144 7694 9178
rect 7518 8886 7694 8920
rect 7518 8628 7694 8662
rect 18175 10318 18209 10654
rect 21833 10318 21867 10654
rect 25491 10318 25525 10654
rect 18175 9830 18209 10166
rect 21833 9830 21867 10166
rect 25491 9830 25525 10166
rect 7518 7899 7694 7933
rect 7518 7441 7694 7475
rect 7518 6609 7694 6643
rect 7518 6151 7694 6185
rect 7518 5319 7694 5353
rect 7518 4861 7694 4895
rect 7518 4029 7694 4063
rect 7518 3571 7694 3605
rect 7518 3448 7694 3482
rect 7518 2990 7694 3024
<< psubdiff >>
rect 4640 28750 4700 28784
rect 10001 28750 10061 28784
rect 4640 28724 4674 28750
rect 3363 27135 3459 27169
rect 4215 27135 4311 27169
rect 3363 27073 3397 27135
rect 4277 27073 4311 27135
rect 3363 25883 3397 25945
rect 4277 25883 4311 25945
rect 3363 25849 3459 25883
rect 4215 25849 4311 25883
rect 10027 28724 10061 28750
rect 4640 25356 4674 25382
rect 10027 25356 10061 25382
rect 4640 25322 4700 25356
rect 10001 25322 10061 25356
rect 22135 25277 22195 25311
rect 24177 25277 24237 25311
rect 22135 25251 22169 25277
rect 11926 24855 11986 24889
rect 20155 24855 20215 24889
rect 11926 24829 11960 24855
rect 20181 24829 20215 24855
rect 11926 23580 11960 23606
rect 20181 23580 20215 23606
rect 11926 23546 11986 23580
rect 20155 23546 20215 23580
rect 24203 25251 24237 25277
rect 22135 23107 22169 23133
rect 25311 24112 25371 24146
rect 25970 24112 26030 24146
rect 25311 24086 25345 24112
rect 25996 24086 26030 24112
rect 25311 23620 25345 23646
rect 25996 23620 26030 23646
rect 25311 23586 25371 23620
rect 25970 23586 26030 23620
rect 24203 23107 24237 23133
rect 22135 23073 22195 23107
rect 24177 23073 24237 23107
rect 24759 23112 24855 23146
rect 25995 23112 26091 23146
rect 24759 23050 24793 23112
rect 26057 23050 26091 23112
rect 22480 22830 22576 22864
rect 23832 22830 23928 22864
rect 22480 22768 22514 22830
rect 15838 22508 15898 22542
rect 16480 22508 16540 22542
rect 15838 22482 15872 22508
rect 12190 21680 12250 21714
rect 14959 21680 15019 21714
rect 12190 21654 12224 21680
rect 14985 21654 15019 21680
rect 12190 15172 12224 15198
rect 16506 22482 16540 22508
rect 15838 17048 15872 17074
rect 23894 22768 23928 22830
rect 24759 22850 24793 22912
rect 26057 22850 26091 22912
rect 24759 22816 24855 22850
rect 25995 22816 26091 22850
rect 22480 21920 22514 21982
rect 23894 21920 23928 21982
rect 22480 21886 22576 21920
rect 23832 21886 23928 21920
rect 16506 17048 16540 17074
rect 15838 17014 15898 17048
rect 16480 17014 16540 17048
rect 14985 15172 15019 15198
rect 12190 15138 12250 15172
rect 14959 15138 15019 15172
rect 15236 16359 16524 16392
rect 15236 16325 15294 16359
rect 15328 16325 15384 16359
rect 15418 16325 15474 16359
rect 15508 16325 15564 16359
rect 15598 16325 15654 16359
rect 15688 16325 15744 16359
rect 15778 16325 15834 16359
rect 15868 16325 15924 16359
rect 15958 16325 16014 16359
rect 16048 16325 16104 16359
rect 16138 16325 16194 16359
rect 16228 16325 16284 16359
rect 16318 16325 16374 16359
rect 16408 16325 16524 16359
rect 15236 16291 16524 16325
rect 15236 16258 15337 16291
rect 15236 16224 15271 16258
rect 15305 16224 15337 16258
rect 16423 16258 16524 16291
rect 15236 16168 15337 16224
rect 15236 16134 15271 16168
rect 15305 16134 15337 16168
rect 15236 16078 15337 16134
rect 15236 16044 15271 16078
rect 15305 16044 15337 16078
rect 15236 15988 15337 16044
rect 15236 15954 15271 15988
rect 15305 15954 15337 15988
rect 15236 15898 15337 15954
rect 15236 15864 15271 15898
rect 15305 15864 15337 15898
rect 15236 15808 15337 15864
rect 15236 15774 15271 15808
rect 15305 15774 15337 15808
rect 15236 15718 15337 15774
rect 15236 15684 15271 15718
rect 15305 15684 15337 15718
rect 15236 15628 15337 15684
rect 15236 15594 15271 15628
rect 15305 15594 15337 15628
rect 15236 15538 15337 15594
rect 15236 15504 15271 15538
rect 15305 15504 15337 15538
rect 15236 15448 15337 15504
rect 15236 15414 15271 15448
rect 15305 15414 15337 15448
rect 15236 15358 15337 15414
rect 15236 15324 15271 15358
rect 15305 15324 15337 15358
rect 15236 15268 15337 15324
rect 15236 15234 15271 15268
rect 15305 15234 15337 15268
rect 16423 16224 16458 16258
rect 16492 16224 16524 16258
rect 16423 16168 16524 16224
rect 16423 16134 16458 16168
rect 16492 16134 16524 16168
rect 16423 16078 16524 16134
rect 16423 16044 16458 16078
rect 16492 16044 16524 16078
rect 16423 15988 16524 16044
rect 16423 15954 16458 15988
rect 16492 15954 16524 15988
rect 16423 15898 16524 15954
rect 16423 15864 16458 15898
rect 16492 15864 16524 15898
rect 16423 15808 16524 15864
rect 16423 15774 16458 15808
rect 16492 15774 16524 15808
rect 16423 15718 16524 15774
rect 16423 15684 16458 15718
rect 16492 15684 16524 15718
rect 16423 15628 16524 15684
rect 16423 15594 16458 15628
rect 16492 15594 16524 15628
rect 16423 15538 16524 15594
rect 16423 15504 16458 15538
rect 16492 15504 16524 15538
rect 16423 15448 16524 15504
rect 16423 15414 16458 15448
rect 16492 15414 16524 15448
rect 16423 15358 16524 15414
rect 16423 15324 16458 15358
rect 16492 15324 16524 15358
rect 16423 15268 16524 15324
rect 15236 15205 15337 15234
rect 16423 15234 16458 15268
rect 16492 15234 16524 15268
rect 16423 15205 16524 15234
rect 15236 15172 16524 15205
rect 15236 15138 15294 15172
rect 15328 15138 15384 15172
rect 15418 15138 15474 15172
rect 15508 15138 15564 15172
rect 15598 15138 15654 15172
rect 15688 15138 15744 15172
rect 15778 15138 15834 15172
rect 15868 15138 15924 15172
rect 15958 15138 16014 15172
rect 16048 15138 16104 15172
rect 16138 15138 16194 15172
rect 16228 15138 16284 15172
rect 16318 15138 16374 15172
rect 16408 15138 16524 15172
rect 15236 15104 16524 15138
rect 5871 10391 7159 10425
rect 2825 10357 2885 10391
rect 5594 10357 5654 10391
rect 2825 10331 2859 10357
rect 5620 10331 5654 10357
rect 2825 3849 2859 3875
rect 5871 10357 5929 10391
rect 5963 10357 6019 10391
rect 6053 10357 6109 10391
rect 6143 10357 6199 10391
rect 6233 10357 6289 10391
rect 6323 10357 6379 10391
rect 6413 10357 6469 10391
rect 6503 10357 6559 10391
rect 6593 10357 6649 10391
rect 6683 10357 6739 10391
rect 6773 10357 6829 10391
rect 6863 10357 6919 10391
rect 6953 10357 7009 10391
rect 7043 10357 7159 10391
rect 5871 10324 7159 10357
rect 5871 10295 5972 10324
rect 5871 10261 5906 10295
rect 5940 10261 5972 10295
rect 7058 10295 7159 10324
rect 5871 10205 5972 10261
rect 5871 10171 5906 10205
rect 5940 10171 5972 10205
rect 5871 10115 5972 10171
rect 5871 10081 5906 10115
rect 5940 10081 5972 10115
rect 5871 10025 5972 10081
rect 5871 9991 5906 10025
rect 5940 9991 5972 10025
rect 5871 9935 5972 9991
rect 5871 9901 5906 9935
rect 5940 9901 5972 9935
rect 5871 9845 5972 9901
rect 5871 9811 5906 9845
rect 5940 9811 5972 9845
rect 5871 9755 5972 9811
rect 5871 9721 5906 9755
rect 5940 9721 5972 9755
rect 5871 9665 5972 9721
rect 5871 9631 5906 9665
rect 5940 9631 5972 9665
rect 5871 9575 5972 9631
rect 5871 9541 5906 9575
rect 5940 9541 5972 9575
rect 5871 9485 5972 9541
rect 5871 9451 5906 9485
rect 5940 9451 5972 9485
rect 5871 9395 5972 9451
rect 5871 9361 5906 9395
rect 5940 9361 5972 9395
rect 5871 9305 5972 9361
rect 5871 9271 5906 9305
rect 5940 9271 5972 9305
rect 7058 10261 7093 10295
rect 7127 10261 7159 10295
rect 7058 10205 7159 10261
rect 7058 10171 7093 10205
rect 7127 10171 7159 10205
rect 7058 10115 7159 10171
rect 7058 10081 7093 10115
rect 7127 10081 7159 10115
rect 7058 10025 7159 10081
rect 7058 9991 7093 10025
rect 7127 9991 7159 10025
rect 7058 9935 7159 9991
rect 7058 9901 7093 9935
rect 7127 9901 7159 9935
rect 7058 9845 7159 9901
rect 7058 9811 7093 9845
rect 7127 9811 7159 9845
rect 7058 9755 7159 9811
rect 7058 9721 7093 9755
rect 7127 9721 7159 9755
rect 7058 9665 7159 9721
rect 7058 9631 7093 9665
rect 7127 9631 7159 9665
rect 7058 9575 7159 9631
rect 7058 9541 7093 9575
rect 7127 9541 7159 9575
rect 7058 9485 7159 9541
rect 7058 9451 7093 9485
rect 7127 9451 7159 9485
rect 7058 9395 7159 9451
rect 7058 9361 7093 9395
rect 7127 9361 7159 9395
rect 7058 9305 7159 9361
rect 5871 9238 5972 9271
rect 7058 9271 7093 9305
rect 7127 9271 7159 9305
rect 7058 9238 7159 9271
rect 5871 9204 7159 9238
rect 5871 9170 5929 9204
rect 5963 9170 6019 9204
rect 6053 9170 6109 9204
rect 6143 9170 6199 9204
rect 6233 9170 6289 9204
rect 6323 9170 6379 9204
rect 6413 9170 6469 9204
rect 6503 9170 6559 9204
rect 6593 9170 6649 9204
rect 6683 9170 6739 9204
rect 6773 9170 6829 9204
rect 6863 9170 6919 9204
rect 6953 9170 7009 9204
rect 7043 9170 7159 9204
rect 5871 9137 7159 9170
rect 19149 8964 19209 8998
rect 24510 8964 24570 8998
rect 19149 8938 19183 8964
rect 5620 3849 5654 3875
rect 2825 3815 2885 3849
rect 5594 3815 5654 3849
rect 6473 8382 6533 8416
rect 7115 8382 7175 8416
rect 6473 8356 6507 8382
rect 7141 8356 7175 8382
rect 6473 2922 6507 2948
rect 17872 7349 17968 7383
rect 18724 7349 18820 7383
rect 17872 7287 17906 7349
rect 18786 7287 18820 7349
rect 17872 6097 17906 6159
rect 18786 6097 18820 6159
rect 17872 6063 17968 6097
rect 18724 6063 18820 6097
rect 24536 8938 24570 8964
rect 19149 5570 19183 5596
rect 24536 5570 24570 5596
rect 19149 5536 19209 5570
rect 24510 5536 24570 5570
rect 7141 2922 7175 2948
rect 6473 2888 6533 2922
rect 7115 2888 7175 2922
<< nsubdiff >>
rect 11874 32908 11934 32942
rect 14214 32908 14274 32942
rect 11874 32882 11908 32908
rect 3409 30711 3469 30745
rect 11157 30711 11217 30745
rect 3409 30685 3443 30711
rect 11183 30685 11217 30711
rect 3409 29403 3443 29429
rect 11183 29403 11217 29429
rect 3409 29369 3469 29403
rect 11157 29369 11217 29403
rect 14240 32882 14274 32908
rect 11874 25321 11908 25347
rect 20795 27824 20855 27858
rect 25541 27824 25601 27858
rect 20795 27798 20829 27824
rect 16853 27146 16949 27180
rect 18691 27146 18787 27180
rect 16853 27084 16887 27146
rect 18753 27084 18787 27146
rect 16853 25448 16887 25510
rect 25567 27798 25601 27824
rect 20795 25559 20829 25585
rect 25567 25559 25601 25585
rect 20795 25525 20855 25559
rect 25541 25525 25601 25559
rect 18753 25448 18787 25510
rect 16853 25414 16949 25448
rect 18691 25414 18787 25448
rect 14240 25321 14274 25347
rect 11874 25287 11934 25321
rect 14214 25287 14274 25321
rect 25279 25126 25375 25160
rect 25573 25126 25731 25160
rect 25929 25126 26025 25160
rect 25279 25064 25313 25126
rect 25635 25064 25669 25126
rect 25279 24308 25313 24370
rect 25991 25064 26025 25126
rect 25635 24308 25669 24370
rect 25991 24308 26025 24370
rect 25279 24274 25375 24308
rect 25573 24274 25731 24308
rect 25929 24274 26025 24308
rect 16712 22516 16772 22550
rect 17196 22516 17256 22550
rect 16712 22490 16746 22516
rect 17222 22490 17256 22516
rect 16712 21300 16746 21326
rect 17222 21300 17256 21326
rect 16712 21266 16772 21300
rect 17196 21266 17256 21300
rect 16688 20649 16784 20683
rect 17158 20649 17254 20683
rect 16688 20587 16722 20649
rect 17220 20587 17254 20649
rect 16688 19997 16722 20059
rect 17220 19997 17254 20059
rect 16688 19963 16784 19997
rect 17158 19963 17254 19997
rect 16688 19359 16784 19393
rect 17158 19359 17254 19393
rect 16688 19297 16722 19359
rect 17220 19297 17254 19359
rect 16688 18707 16722 18769
rect 17220 18707 17254 18769
rect 16688 18673 16784 18707
rect 17158 18673 17254 18707
rect 16688 18069 16784 18103
rect 17158 18069 17254 18103
rect 16688 18007 16722 18069
rect 17220 18007 17254 18069
rect 16688 17417 16722 17479
rect 17220 17417 17254 17479
rect 16688 17383 16784 17417
rect 17158 17383 17254 17417
rect 16697 16968 16780 17017
rect 17159 16968 17247 17017
rect 16697 16906 16745 16968
rect 17195 16899 17247 16968
rect 15399 16210 16361 16229
rect 15399 16176 15494 16210
rect 15528 16176 15584 16210
rect 15618 16176 15674 16210
rect 15708 16176 15764 16210
rect 15798 16176 15854 16210
rect 15888 16176 15944 16210
rect 15978 16176 16034 16210
rect 16068 16176 16124 16210
rect 16158 16176 16214 16210
rect 16248 16176 16361 16210
rect 15399 16157 16361 16176
rect 15399 16152 15471 16157
rect 15399 16118 15418 16152
rect 15452 16118 15471 16152
rect 15399 16062 15471 16118
rect 16289 16118 16361 16157
rect 15399 16028 15418 16062
rect 15452 16028 15471 16062
rect 15399 15972 15471 16028
rect 15399 15938 15418 15972
rect 15452 15938 15471 15972
rect 15399 15882 15471 15938
rect 15399 15848 15418 15882
rect 15452 15848 15471 15882
rect 15399 15792 15471 15848
rect 15399 15758 15418 15792
rect 15452 15758 15471 15792
rect 15399 15702 15471 15758
rect 15399 15668 15418 15702
rect 15452 15668 15471 15702
rect 15399 15612 15471 15668
rect 15399 15578 15418 15612
rect 15452 15578 15471 15612
rect 15399 15522 15471 15578
rect 15399 15488 15418 15522
rect 15452 15488 15471 15522
rect 15399 15432 15471 15488
rect 15399 15398 15418 15432
rect 15452 15398 15471 15432
rect 16289 16084 16308 16118
rect 16342 16084 16361 16118
rect 16289 16028 16361 16084
rect 16289 15994 16308 16028
rect 16342 15994 16361 16028
rect 16289 15938 16361 15994
rect 16289 15904 16308 15938
rect 16342 15904 16361 15938
rect 16289 15848 16361 15904
rect 16289 15814 16308 15848
rect 16342 15814 16361 15848
rect 16289 15758 16361 15814
rect 16289 15724 16308 15758
rect 16342 15724 16361 15758
rect 16289 15668 16361 15724
rect 16289 15634 16308 15668
rect 16342 15634 16361 15668
rect 16289 15578 16361 15634
rect 16289 15544 16308 15578
rect 16342 15544 16361 15578
rect 16289 15488 16361 15544
rect 16289 15454 16308 15488
rect 16342 15454 16361 15488
rect 15399 15339 15471 15398
rect 16289 15398 16361 15454
rect 16289 15364 16308 15398
rect 16342 15364 16361 15398
rect 16289 15339 16361 15364
rect 15399 15320 16361 15339
rect 15399 15286 15475 15320
rect 15509 15286 15565 15320
rect 15599 15286 15655 15320
rect 15689 15286 15745 15320
rect 15779 15286 15835 15320
rect 15869 15286 15925 15320
rect 15959 15286 16015 15320
rect 16049 15286 16105 15320
rect 16139 15286 16195 15320
rect 16229 15286 16361 15320
rect 15399 15267 16361 15286
rect 16697 16372 16745 16629
rect 16697 15128 16745 15264
rect 17195 15128 17247 15224
rect 16697 15076 16864 15128
rect 17100 15076 17247 15128
rect 17918 10925 17978 10959
rect 25666 10925 25726 10959
rect 17918 10899 17952 10925
rect 6034 10243 6996 10262
rect 6034 10209 6110 10243
rect 6144 10209 6200 10243
rect 6234 10209 6290 10243
rect 6324 10209 6380 10243
rect 6414 10209 6470 10243
rect 6504 10209 6560 10243
rect 6594 10209 6650 10243
rect 6684 10209 6740 10243
rect 6774 10209 6830 10243
rect 6864 10209 6996 10243
rect 6034 10190 6996 10209
rect 6034 10131 6106 10190
rect 6034 10097 6053 10131
rect 6087 10097 6106 10131
rect 6924 10165 6996 10190
rect 6924 10131 6943 10165
rect 6977 10131 6996 10165
rect 6034 10041 6106 10097
rect 6034 10007 6053 10041
rect 6087 10007 6106 10041
rect 6034 9951 6106 10007
rect 6034 9917 6053 9951
rect 6087 9917 6106 9951
rect 6034 9861 6106 9917
rect 6034 9827 6053 9861
rect 6087 9827 6106 9861
rect 6034 9771 6106 9827
rect 6034 9737 6053 9771
rect 6087 9737 6106 9771
rect 6034 9681 6106 9737
rect 6034 9647 6053 9681
rect 6087 9647 6106 9681
rect 6034 9591 6106 9647
rect 6034 9557 6053 9591
rect 6087 9557 6106 9591
rect 6034 9501 6106 9557
rect 6034 9467 6053 9501
rect 6087 9467 6106 9501
rect 6034 9411 6106 9467
rect 6924 10075 6996 10131
rect 6924 10041 6943 10075
rect 6977 10041 6996 10075
rect 6924 9985 6996 10041
rect 6924 9951 6943 9985
rect 6977 9951 6996 9985
rect 6924 9895 6996 9951
rect 6924 9861 6943 9895
rect 6977 9861 6996 9895
rect 6924 9805 6996 9861
rect 6924 9771 6943 9805
rect 6977 9771 6996 9805
rect 6924 9715 6996 9771
rect 6924 9681 6943 9715
rect 6977 9681 6996 9715
rect 6924 9625 6996 9681
rect 6924 9591 6943 9625
rect 6977 9591 6996 9625
rect 6924 9535 6996 9591
rect 6924 9501 6943 9535
rect 6977 9501 6996 9535
rect 6924 9445 6996 9501
rect 6034 9377 6053 9411
rect 6087 9377 6106 9411
rect 6034 9372 6106 9377
rect 6924 9411 6943 9445
rect 6977 9411 6996 9445
rect 6924 9372 6996 9411
rect 6034 9353 6996 9372
rect 6034 9319 6129 9353
rect 6163 9319 6219 9353
rect 6253 9319 6309 9353
rect 6343 9319 6399 9353
rect 6433 9319 6489 9353
rect 6523 9319 6579 9353
rect 6613 9319 6669 9353
rect 6703 9319 6759 9353
rect 6793 9319 6849 9353
rect 6883 9319 6996 9353
rect 6034 9300 6996 9319
rect 7332 10401 7499 10453
rect 7735 10401 7882 10453
rect 7332 10265 7380 10401
rect 7830 10305 7882 10401
rect 7332 8900 7380 9157
rect 7332 8561 7380 8623
rect 25692 10899 25726 10925
rect 17918 9617 17952 9643
rect 25692 9617 25726 9643
rect 17918 9583 17978 9617
rect 25666 9583 25726 9617
rect 7830 8561 7882 8630
rect 7332 8512 7415 8561
rect 7794 8512 7882 8561
rect 7323 8013 7419 8047
rect 7793 8013 7889 8047
rect 7323 7951 7357 8013
rect 7855 7951 7889 8013
rect 7323 7361 7357 7423
rect 7855 7361 7889 7423
rect 7323 7327 7419 7361
rect 7793 7327 7889 7361
rect 7323 6723 7419 6757
rect 7793 6723 7889 6757
rect 7323 6661 7357 6723
rect 7855 6661 7889 6723
rect 7323 6071 7357 6133
rect 7855 6071 7889 6133
rect 7323 6037 7419 6071
rect 7793 6037 7889 6071
rect 7323 5433 7419 5467
rect 7793 5433 7889 5467
rect 7323 5371 7357 5433
rect 7855 5371 7889 5433
rect 7323 4781 7357 4843
rect 7855 4781 7889 4843
rect 7323 4747 7419 4781
rect 7793 4747 7889 4781
rect 7347 4130 7407 4164
rect 7831 4130 7891 4164
rect 7347 4104 7381 4130
rect 7857 4104 7891 4130
rect 7347 2914 7381 2940
rect 7857 2914 7891 2940
rect 7347 2880 7407 2914
rect 7831 2880 7891 2914
<< psubdiffcont >>
rect 4700 28750 10001 28784
rect 3459 27135 4215 27169
rect 3363 25945 3397 27073
rect 4277 25945 4311 27073
rect 3459 25849 4215 25883
rect 4640 25382 4674 28724
rect 10027 25382 10061 28724
rect 4700 25322 10001 25356
rect 22195 25277 24177 25311
rect 11986 24855 20155 24889
rect 11926 23606 11960 24829
rect 20181 23606 20215 24829
rect 11986 23546 20155 23580
rect 22135 23133 22169 25251
rect 24203 23133 24237 25251
rect 25371 24112 25970 24146
rect 25311 23646 25345 24086
rect 25996 23646 26030 24086
rect 25371 23586 25970 23620
rect 22195 23073 24177 23107
rect 24855 23112 25995 23146
rect 24759 22912 24793 23050
rect 22576 22830 23832 22864
rect 15898 22508 16480 22542
rect 12250 21680 14959 21714
rect 12190 15198 12224 21654
rect 14985 15198 15019 21654
rect 15838 17074 15872 22482
rect 16506 17074 16540 22482
rect 22480 21982 22514 22768
rect 26057 22912 26091 23050
rect 24855 22816 25995 22850
rect 23894 21982 23928 22768
rect 22576 21886 23832 21920
rect 15898 17014 16480 17048
rect 12250 15138 14959 15172
rect 15294 16325 15328 16359
rect 15384 16325 15418 16359
rect 15474 16325 15508 16359
rect 15564 16325 15598 16359
rect 15654 16325 15688 16359
rect 15744 16325 15778 16359
rect 15834 16325 15868 16359
rect 15924 16325 15958 16359
rect 16014 16325 16048 16359
rect 16104 16325 16138 16359
rect 16194 16325 16228 16359
rect 16284 16325 16318 16359
rect 16374 16325 16408 16359
rect 15271 16224 15305 16258
rect 15271 16134 15305 16168
rect 15271 16044 15305 16078
rect 15271 15954 15305 15988
rect 15271 15864 15305 15898
rect 15271 15774 15305 15808
rect 15271 15684 15305 15718
rect 15271 15594 15305 15628
rect 15271 15504 15305 15538
rect 15271 15414 15305 15448
rect 15271 15324 15305 15358
rect 15271 15234 15305 15268
rect 16458 16224 16492 16258
rect 16458 16134 16492 16168
rect 16458 16044 16492 16078
rect 16458 15954 16492 15988
rect 16458 15864 16492 15898
rect 16458 15774 16492 15808
rect 16458 15684 16492 15718
rect 16458 15594 16492 15628
rect 16458 15504 16492 15538
rect 16458 15414 16492 15448
rect 16458 15324 16492 15358
rect 16458 15234 16492 15268
rect 15294 15138 15328 15172
rect 15384 15138 15418 15172
rect 15474 15138 15508 15172
rect 15564 15138 15598 15172
rect 15654 15138 15688 15172
rect 15744 15138 15778 15172
rect 15834 15138 15868 15172
rect 15924 15138 15958 15172
rect 16014 15138 16048 15172
rect 16104 15138 16138 15172
rect 16194 15138 16228 15172
rect 16284 15138 16318 15172
rect 16374 15138 16408 15172
rect 2885 10357 5594 10391
rect 2825 3875 2859 10331
rect 5620 3875 5654 10331
rect 5929 10357 5963 10391
rect 6019 10357 6053 10391
rect 6109 10357 6143 10391
rect 6199 10357 6233 10391
rect 6289 10357 6323 10391
rect 6379 10357 6413 10391
rect 6469 10357 6503 10391
rect 6559 10357 6593 10391
rect 6649 10357 6683 10391
rect 6739 10357 6773 10391
rect 6829 10357 6863 10391
rect 6919 10357 6953 10391
rect 7009 10357 7043 10391
rect 5906 10261 5940 10295
rect 5906 10171 5940 10205
rect 5906 10081 5940 10115
rect 5906 9991 5940 10025
rect 5906 9901 5940 9935
rect 5906 9811 5940 9845
rect 5906 9721 5940 9755
rect 5906 9631 5940 9665
rect 5906 9541 5940 9575
rect 5906 9451 5940 9485
rect 5906 9361 5940 9395
rect 5906 9271 5940 9305
rect 7093 10261 7127 10295
rect 7093 10171 7127 10205
rect 7093 10081 7127 10115
rect 7093 9991 7127 10025
rect 7093 9901 7127 9935
rect 7093 9811 7127 9845
rect 7093 9721 7127 9755
rect 7093 9631 7127 9665
rect 7093 9541 7127 9575
rect 7093 9451 7127 9485
rect 7093 9361 7127 9395
rect 7093 9271 7127 9305
rect 5929 9170 5963 9204
rect 6019 9170 6053 9204
rect 6109 9170 6143 9204
rect 6199 9170 6233 9204
rect 6289 9170 6323 9204
rect 6379 9170 6413 9204
rect 6469 9170 6503 9204
rect 6559 9170 6593 9204
rect 6649 9170 6683 9204
rect 6739 9170 6773 9204
rect 6829 9170 6863 9204
rect 6919 9170 6953 9204
rect 7009 9170 7043 9204
rect 19209 8964 24510 8998
rect 2885 3815 5594 3849
rect 6533 8382 7115 8416
rect 6473 2948 6507 8356
rect 7141 2948 7175 8356
rect 17968 7349 18724 7383
rect 17872 6159 17906 7287
rect 18786 6159 18820 7287
rect 17968 6063 18724 6097
rect 19149 5596 19183 8938
rect 24536 5596 24570 8938
rect 19209 5536 24510 5570
rect 6533 2888 7115 2922
<< nsubdiffcont >>
rect 11934 32908 14214 32942
rect 3469 30711 11157 30745
rect 3409 29429 3443 30685
rect 11183 29429 11217 30685
rect 3469 29369 11157 29403
rect 11874 25347 11908 32882
rect 14240 25347 14274 32882
rect 20855 27824 25541 27858
rect 16949 27146 18691 27180
rect 16853 25510 16887 27084
rect 18753 25510 18787 27084
rect 20795 25585 20829 27798
rect 25567 25585 25601 27798
rect 20855 25525 25541 25559
rect 16949 25414 18691 25448
rect 11934 25287 14214 25321
rect 25375 25126 25573 25160
rect 25731 25126 25929 25160
rect 25279 24370 25313 25064
rect 25635 24370 25669 25064
rect 25991 24370 26025 25064
rect 25375 24274 25573 24308
rect 25731 24274 25929 24308
rect 16772 22516 17196 22550
rect 16712 21326 16746 22490
rect 17222 21326 17256 22490
rect 16772 21266 17196 21300
rect 16784 20649 17158 20683
rect 16688 20059 16722 20587
rect 17220 20059 17254 20587
rect 16784 19963 17158 19997
rect 16784 19359 17158 19393
rect 16688 18769 16722 19297
rect 17220 18769 17254 19297
rect 16784 18673 17158 18707
rect 16784 18069 17158 18103
rect 16688 17479 16722 18007
rect 17220 17479 17254 18007
rect 16784 17383 17158 17417
rect 16780 16968 17159 17017
rect 16697 16629 16745 16906
rect 15494 16176 15528 16210
rect 15584 16176 15618 16210
rect 15674 16176 15708 16210
rect 15764 16176 15798 16210
rect 15854 16176 15888 16210
rect 15944 16176 15978 16210
rect 16034 16176 16068 16210
rect 16124 16176 16158 16210
rect 16214 16176 16248 16210
rect 15418 16118 15452 16152
rect 15418 16028 15452 16062
rect 15418 15938 15452 15972
rect 15418 15848 15452 15882
rect 15418 15758 15452 15792
rect 15418 15668 15452 15702
rect 15418 15578 15452 15612
rect 15418 15488 15452 15522
rect 15418 15398 15452 15432
rect 16308 16084 16342 16118
rect 16308 15994 16342 16028
rect 16308 15904 16342 15938
rect 16308 15814 16342 15848
rect 16308 15724 16342 15758
rect 16308 15634 16342 15668
rect 16308 15544 16342 15578
rect 16308 15454 16342 15488
rect 16308 15364 16342 15398
rect 15475 15286 15509 15320
rect 15565 15286 15599 15320
rect 15655 15286 15689 15320
rect 15745 15286 15779 15320
rect 15835 15286 15869 15320
rect 15925 15286 15959 15320
rect 16015 15286 16049 15320
rect 16105 15286 16139 15320
rect 16195 15286 16229 15320
rect 16697 15264 16745 16372
rect 17195 15224 17247 16899
rect 16864 15076 17100 15128
rect 17978 10925 25666 10959
rect 6110 10209 6144 10243
rect 6200 10209 6234 10243
rect 6290 10209 6324 10243
rect 6380 10209 6414 10243
rect 6470 10209 6504 10243
rect 6560 10209 6594 10243
rect 6650 10209 6684 10243
rect 6740 10209 6774 10243
rect 6830 10209 6864 10243
rect 6053 10097 6087 10131
rect 6943 10131 6977 10165
rect 6053 10007 6087 10041
rect 6053 9917 6087 9951
rect 6053 9827 6087 9861
rect 6053 9737 6087 9771
rect 6053 9647 6087 9681
rect 6053 9557 6087 9591
rect 6053 9467 6087 9501
rect 6943 10041 6977 10075
rect 6943 9951 6977 9985
rect 6943 9861 6977 9895
rect 6943 9771 6977 9805
rect 6943 9681 6977 9715
rect 6943 9591 6977 9625
rect 6943 9501 6977 9535
rect 6053 9377 6087 9411
rect 6943 9411 6977 9445
rect 6129 9319 6163 9353
rect 6219 9319 6253 9353
rect 6309 9319 6343 9353
rect 6399 9319 6433 9353
rect 6489 9319 6523 9353
rect 6579 9319 6613 9353
rect 6669 9319 6703 9353
rect 6759 9319 6793 9353
rect 6849 9319 6883 9353
rect 7499 10401 7735 10453
rect 7332 9157 7380 10265
rect 7332 8623 7380 8900
rect 7830 8630 7882 10305
rect 17918 9643 17952 10899
rect 25692 9643 25726 10899
rect 17978 9583 25666 9617
rect 7415 8512 7794 8561
rect 7419 8013 7793 8047
rect 7323 7423 7357 7951
rect 7855 7423 7889 7951
rect 7419 7327 7793 7361
rect 7419 6723 7793 6757
rect 7323 6133 7357 6661
rect 7855 6133 7889 6661
rect 7419 6037 7793 6071
rect 7419 5433 7793 5467
rect 7323 4843 7357 5371
rect 7855 4843 7889 5371
rect 7419 4747 7793 4781
rect 7407 4130 7831 4164
rect 7347 2940 7381 4104
rect 7857 2940 7891 4104
rect 7407 2880 7831 2914
<< poly >>
rect 3712 30533 7312 30549
rect 3712 30499 3728 30533
rect 7296 30499 7312 30533
rect 3712 30452 7312 30499
rect 7370 30533 10970 30549
rect 7370 30499 7386 30533
rect 10954 30499 10970 30533
rect 7370 30452 10970 30499
rect 3712 30045 7312 30092
rect 3712 30011 3728 30045
rect 7296 30011 7312 30045
rect 3712 29964 7312 30011
rect 7370 30045 10970 30092
rect 7370 30011 7386 30045
rect 10954 30011 10970 30045
rect 7370 29964 10970 30011
rect 3712 29557 7312 29604
rect 3712 29523 3728 29557
rect 7296 29523 7312 29557
rect 3712 29507 7312 29523
rect 7370 29557 10970 29604
rect 7370 29523 7386 29557
rect 10954 29523 10970 29557
rect 7370 29507 10970 29523
rect 3449 26993 3537 27009
rect 3449 26025 3465 26993
rect 3499 26025 3537 26993
rect 3449 26009 3537 26025
rect 4137 26993 4225 27009
rect 4137 26025 4175 26993
rect 4209 26025 4225 26993
rect 4137 26009 4225 26025
rect 4922 28652 7322 28668
rect 4922 28618 4938 28652
rect 7306 28618 7322 28652
rect 4922 28580 7322 28618
rect 7380 28652 9780 28668
rect 7380 28618 7396 28652
rect 9764 28618 9780 28652
rect 7380 28580 9780 28618
rect 4922 27342 7322 27380
rect 4922 27308 4938 27342
rect 7306 27308 7322 27342
rect 4922 27292 7322 27308
rect 7380 27342 9780 27380
rect 7380 27308 7396 27342
rect 9764 27308 9780 27342
rect 7380 27292 9780 27308
rect 4921 26777 7321 26793
rect 4921 26743 4937 26777
rect 7305 26743 7321 26777
rect 4921 26705 7321 26743
rect 7379 26777 9779 26793
rect 7379 26743 7395 26777
rect 9763 26743 9779 26777
rect 7379 26705 9779 26743
rect 4921 25467 7321 25505
rect 4921 25433 4937 25467
rect 7305 25433 7321 25467
rect 4921 25417 7321 25433
rect 7379 25467 9779 25505
rect 7379 25433 7395 25467
rect 9763 25433 9779 25467
rect 7379 25417 9779 25433
rect 12184 32609 12564 32625
rect 12184 32575 12200 32609
rect 12548 32575 12564 32609
rect 12184 32528 12564 32575
rect 12622 32609 13002 32625
rect 12622 32575 12638 32609
rect 12986 32575 13002 32609
rect 12622 32528 13002 32575
rect 13060 32609 13440 32625
rect 13060 32575 13076 32609
rect 13424 32575 13440 32609
rect 13060 32528 13440 32575
rect 13498 32609 13878 32625
rect 13498 32575 13514 32609
rect 13862 32575 13878 32609
rect 13498 32528 13878 32575
rect 12184 29481 12564 29528
rect 12184 29447 12200 29481
rect 12548 29447 12564 29481
rect 12184 29431 12564 29447
rect 12622 29481 13002 29528
rect 12622 29447 12638 29481
rect 12986 29447 13002 29481
rect 12622 29431 13002 29447
rect 13060 29481 13440 29528
rect 13060 29447 13076 29481
rect 13424 29447 13440 29481
rect 13060 29431 13440 29447
rect 13498 29481 13878 29528
rect 13498 29447 13514 29481
rect 13862 29447 13878 29481
rect 13498 29431 13878 29447
rect 12184 28632 12564 28648
rect 12184 28598 12200 28632
rect 12548 28598 12564 28632
rect 12184 28551 12564 28598
rect 12622 28632 13002 28648
rect 12622 28598 12638 28632
rect 12986 28598 13002 28632
rect 12622 28551 13002 28598
rect 13060 28632 13440 28648
rect 13060 28598 13076 28632
rect 13424 28598 13440 28632
rect 13060 28551 13440 28598
rect 13498 28632 13878 28648
rect 13498 28598 13514 28632
rect 13862 28598 13878 28632
rect 13498 28551 13878 28598
rect 12184 25504 12564 25551
rect 12184 25470 12200 25504
rect 12548 25470 12564 25504
rect 12184 25454 12564 25470
rect 12622 25504 13002 25551
rect 12622 25470 12638 25504
rect 12986 25470 13002 25504
rect 12622 25454 13002 25470
rect 13060 25504 13440 25551
rect 13060 25470 13076 25504
rect 13424 25470 13440 25504
rect 13060 25454 13440 25470
rect 13498 25504 13878 25551
rect 13498 25470 13514 25504
rect 13862 25470 13878 25504
rect 13498 25454 13878 25470
rect 17013 27078 17373 27094
rect 17013 27044 17029 27078
rect 17357 27044 17373 27078
rect 17013 26997 17373 27044
rect 17431 27078 17791 27094
rect 17431 27044 17447 27078
rect 17775 27044 17791 27078
rect 17431 26997 17791 27044
rect 17849 27078 18209 27094
rect 17849 27044 17865 27078
rect 18193 27044 18209 27078
rect 17849 26997 18209 27044
rect 18267 27078 18627 27094
rect 18267 27044 18283 27078
rect 18611 27044 18627 27078
rect 18267 26997 18627 27044
rect 17013 25550 17373 25597
rect 17013 25516 17029 25550
rect 17357 25516 17373 25550
rect 17013 25500 17373 25516
rect 17431 25550 17791 25597
rect 17431 25516 17447 25550
rect 17775 25516 17791 25550
rect 17431 25500 17791 25516
rect 17849 25550 18209 25597
rect 17849 25516 17865 25550
rect 18193 25516 18209 25550
rect 17849 25500 18209 25516
rect 18267 25550 18627 25597
rect 18267 25516 18283 25550
rect 18611 25516 18627 25550
rect 18267 25500 18627 25516
rect 21106 27623 22106 27639
rect 21106 27589 21122 27623
rect 22090 27589 22106 27623
rect 21106 27542 22106 27589
rect 22164 27623 23164 27639
rect 22164 27589 22180 27623
rect 23148 27589 23164 27623
rect 22164 27542 23164 27589
rect 23222 27623 24222 27639
rect 23222 27589 23238 27623
rect 24206 27589 24222 27623
rect 23222 27542 24222 27589
rect 24280 27623 25280 27639
rect 24280 27589 24296 27623
rect 25264 27589 25280 27623
rect 24280 27542 25280 27589
rect 21106 26995 22106 27042
rect 21106 26961 21122 26995
rect 22090 26961 22106 26995
rect 21106 26945 22106 26961
rect 22164 26995 23164 27042
rect 22164 26961 22180 26995
rect 23148 26961 23164 26995
rect 22164 26945 23164 26961
rect 23222 26995 24222 27042
rect 23222 26961 23238 26995
rect 24206 26961 24222 26995
rect 23222 26945 24222 26961
rect 24280 26995 25280 27042
rect 24280 26961 24296 26995
rect 25264 26961 25280 26995
rect 24280 26945 25280 26961
rect 21106 26461 22106 26477
rect 21106 26427 21122 26461
rect 22090 26427 22106 26461
rect 21106 26380 22106 26427
rect 22164 26461 23164 26477
rect 22164 26427 22180 26461
rect 23148 26427 23164 26461
rect 22164 26380 23164 26427
rect 23222 26461 24222 26477
rect 23222 26427 23238 26461
rect 24206 26427 24222 26461
rect 23222 26380 24222 26427
rect 24280 26461 25280 26477
rect 24280 26427 24296 26461
rect 25264 26427 25280 26461
rect 24280 26380 25280 26427
rect 21106 25833 22106 25880
rect 21106 25799 21122 25833
rect 22090 25799 22106 25833
rect 21106 25783 22106 25799
rect 22164 25833 23164 25880
rect 22164 25799 22180 25833
rect 23148 25799 23164 25833
rect 22164 25783 23164 25799
rect 23222 25833 24222 25880
rect 23222 25799 23238 25833
rect 24206 25799 24222 25833
rect 23222 25783 24222 25799
rect 24280 25833 25280 25880
rect 24280 25799 24296 25833
rect 25264 25799 25280 25833
rect 24280 25783 25280 25799
rect 12194 24597 14074 24613
rect 12194 24563 12210 24597
rect 14058 24563 14074 24597
rect 12194 24525 14074 24563
rect 14132 24597 16012 24613
rect 14132 24563 14148 24597
rect 15996 24563 16012 24597
rect 14132 24525 16012 24563
rect 16070 24597 17950 24613
rect 16070 24563 16086 24597
rect 17934 24563 17950 24597
rect 16070 24525 17950 24563
rect 18008 24597 19888 24613
rect 18008 24563 18024 24597
rect 19872 24563 19888 24597
rect 18008 24525 19888 24563
rect 12194 24187 14074 24225
rect 12194 24153 12210 24187
rect 14058 24153 14074 24187
rect 12194 24115 14074 24153
rect 14132 24187 16012 24225
rect 14132 24153 14148 24187
rect 15996 24153 16012 24187
rect 14132 24115 16012 24153
rect 16070 24187 17950 24225
rect 16070 24153 16086 24187
rect 17934 24153 17950 24187
rect 16070 24115 17950 24153
rect 18008 24187 19888 24225
rect 18008 24153 18024 24187
rect 19872 24153 19888 24187
rect 18008 24115 19888 24153
rect 12194 23777 14074 23815
rect 12194 23743 12210 23777
rect 14058 23743 14074 23777
rect 12194 23727 14074 23743
rect 14132 23777 16012 23815
rect 14132 23743 14148 23777
rect 15996 23743 16012 23777
rect 14132 23727 16012 23743
rect 16070 23777 17950 23815
rect 16070 23743 16086 23777
rect 17934 23743 17950 23777
rect 16070 23727 17950 23743
rect 18008 23777 19888 23815
rect 18008 23743 18024 23777
rect 19872 23743 19888 23777
rect 18008 23727 19888 23743
rect 22291 25167 22691 25183
rect 22291 25133 22307 25167
rect 22675 25133 22691 25167
rect 22291 25095 22691 25133
rect 22749 25167 23149 25183
rect 22749 25133 22765 25167
rect 23133 25133 23149 25167
rect 22749 25095 23149 25133
rect 23207 25167 23607 25183
rect 23207 25133 23223 25167
rect 23591 25133 23607 25167
rect 23207 25095 23607 25133
rect 23665 25167 24065 25183
rect 23665 25133 23681 25167
rect 24049 25133 24065 25167
rect 23665 25095 24065 25133
rect 22291 24457 22691 24495
rect 22291 24423 22307 24457
rect 22675 24423 22691 24457
rect 22291 24407 22691 24423
rect 22749 24457 23149 24495
rect 22749 24423 22765 24457
rect 23133 24423 23149 24457
rect 22749 24407 23149 24423
rect 23207 24457 23607 24495
rect 23207 24423 23223 24457
rect 23591 24423 23607 24457
rect 23207 24407 23607 24423
rect 23665 24457 24065 24495
rect 23665 24423 23681 24457
rect 24049 24423 24065 24457
rect 23665 24407 24065 24423
rect 22291 23960 22691 23976
rect 22291 23926 22307 23960
rect 22675 23926 22691 23960
rect 22291 23888 22691 23926
rect 22749 23960 23149 23976
rect 22749 23926 22765 23960
rect 23133 23926 23149 23960
rect 22749 23888 23149 23926
rect 23207 23960 23607 23976
rect 23207 23926 23223 23960
rect 23591 23926 23607 23960
rect 23207 23888 23607 23926
rect 23665 23960 24065 23976
rect 23665 23926 23681 23960
rect 24049 23926 24065 23960
rect 23665 23888 24065 23926
rect 22291 23250 22691 23288
rect 22291 23216 22307 23250
rect 22675 23216 22691 23250
rect 22291 23200 22691 23216
rect 22749 23250 23149 23288
rect 22749 23216 22765 23250
rect 23133 23216 23149 23250
rect 22749 23200 23149 23216
rect 23207 23250 23607 23288
rect 23207 23216 23223 23250
rect 23591 23216 23607 23250
rect 23207 23200 23607 23216
rect 23665 23250 24065 23288
rect 23665 23216 23681 23250
rect 24049 23216 24065 23250
rect 23665 23200 24065 23216
rect 25439 25058 25509 25074
rect 25439 25024 25455 25058
rect 25493 25024 25509 25058
rect 25439 24977 25509 25024
rect 25439 24410 25509 24457
rect 25439 24376 25455 24410
rect 25493 24376 25509 24410
rect 25439 24360 25509 24376
rect 25795 25058 25865 25074
rect 25795 25024 25811 25058
rect 25849 25024 25865 25058
rect 25795 24977 25865 25024
rect 25795 24410 25865 24457
rect 25795 24376 25811 24410
rect 25849 24376 25865 24410
rect 25795 24360 25865 24376
rect 25461 24044 25527 24060
rect 25461 24010 25477 24044
rect 25511 24010 25527 24044
rect 25461 23994 25527 24010
rect 25817 24044 25883 24060
rect 25817 24010 25833 24044
rect 25867 24010 25883 24044
rect 25817 23994 25883 24010
rect 25479 23972 25509 23994
rect 25835 23972 25865 23994
rect 25479 23750 25509 23772
rect 25835 23750 25865 23772
rect 25461 23734 25527 23750
rect 25461 23700 25477 23734
rect 25511 23700 25527 23734
rect 25461 23684 25527 23700
rect 25817 23734 25883 23750
rect 25817 23700 25833 23734
rect 25867 23700 25883 23734
rect 25817 23684 25883 23700
rect 12378 21508 12466 21524
rect 12378 21340 12394 21508
rect 12428 21340 12466 21508
rect 12378 21324 12466 21340
rect 13266 21508 13354 21524
rect 13266 21340 13304 21508
rect 13338 21340 13354 21508
rect 13266 21324 13354 21340
rect 13859 21508 13947 21524
rect 13859 21340 13875 21508
rect 13909 21340 13947 21508
rect 13859 21324 13947 21340
rect 14747 21508 14835 21524
rect 14747 21340 14785 21508
rect 14819 21340 14835 21508
rect 14747 21324 14835 21340
rect 12378 21250 12466 21266
rect 12378 21082 12394 21250
rect 12428 21082 12466 21250
rect 12378 21066 12466 21082
rect 13266 21250 13354 21266
rect 13266 21082 13304 21250
rect 13338 21082 13354 21250
rect 13266 21066 13354 21082
rect 13859 21250 13947 21266
rect 13859 21082 13875 21250
rect 13909 21082 13947 21250
rect 13859 21066 13947 21082
rect 14747 21250 14835 21266
rect 14747 21082 14785 21250
rect 14819 21082 14835 21250
rect 14747 21066 14835 21082
rect 12378 20992 12466 21008
rect 12378 20824 12394 20992
rect 12428 20824 12466 20992
rect 12378 20808 12466 20824
rect 13266 20992 13354 21008
rect 13266 20824 13304 20992
rect 13338 20824 13354 20992
rect 13266 20808 13354 20824
rect 13859 20992 13947 21008
rect 13859 20824 13875 20992
rect 13909 20824 13947 20992
rect 13859 20808 13947 20824
rect 14747 20992 14835 21008
rect 14747 20824 14785 20992
rect 14819 20824 14835 20992
rect 14747 20808 14835 20824
rect 12378 20734 12466 20750
rect 12378 20566 12394 20734
rect 12428 20566 12466 20734
rect 12378 20550 12466 20566
rect 13266 20734 13354 20750
rect 13266 20566 13304 20734
rect 13338 20566 13354 20734
rect 13266 20550 13354 20566
rect 13859 20734 13947 20750
rect 13859 20566 13875 20734
rect 13909 20566 13947 20734
rect 13859 20550 13947 20566
rect 14747 20734 14835 20750
rect 14747 20566 14785 20734
rect 14819 20566 14835 20734
rect 14747 20550 14835 20566
rect 12378 20476 12466 20492
rect 12378 20308 12394 20476
rect 12428 20308 12466 20476
rect 12378 20292 12466 20308
rect 13266 20476 13354 20492
rect 13266 20308 13304 20476
rect 13338 20308 13354 20476
rect 13266 20292 13354 20308
rect 13859 20476 13947 20492
rect 13859 20308 13875 20476
rect 13909 20308 13947 20476
rect 13859 20292 13947 20308
rect 14747 20476 14835 20492
rect 14747 20308 14785 20476
rect 14819 20308 14835 20476
rect 14747 20292 14835 20308
rect 12378 20218 12466 20234
rect 12378 20050 12394 20218
rect 12428 20050 12466 20218
rect 12378 20034 12466 20050
rect 13266 20218 13354 20234
rect 13266 20050 13304 20218
rect 13338 20050 13354 20218
rect 13266 20034 13354 20050
rect 13859 20218 13947 20234
rect 13859 20050 13875 20218
rect 13909 20050 13947 20218
rect 13859 20034 13947 20050
rect 14747 20218 14835 20234
rect 14747 20050 14785 20218
rect 14819 20050 14835 20218
rect 14747 20034 14835 20050
rect 12378 19960 12466 19976
rect 12378 19792 12394 19960
rect 12428 19792 12466 19960
rect 12378 19776 12466 19792
rect 13266 19960 13354 19976
rect 13266 19792 13304 19960
rect 13338 19792 13354 19960
rect 13266 19776 13354 19792
rect 13859 19960 13947 19976
rect 13859 19792 13875 19960
rect 13909 19792 13947 19960
rect 13859 19776 13947 19792
rect 14747 19960 14835 19976
rect 14747 19792 14785 19960
rect 14819 19792 14835 19960
rect 14747 19776 14835 19792
rect 12378 19702 12466 19718
rect 12378 19534 12394 19702
rect 12428 19534 12466 19702
rect 12378 19518 12466 19534
rect 13266 19702 13354 19718
rect 13266 19534 13304 19702
rect 13338 19534 13354 19702
rect 13266 19518 13354 19534
rect 13859 19702 13947 19718
rect 13859 19534 13875 19702
rect 13909 19534 13947 19702
rect 13859 19518 13947 19534
rect 14747 19702 14835 19718
rect 14747 19534 14785 19702
rect 14819 19534 14835 19702
rect 14747 19518 14835 19534
rect 12378 19444 12466 19460
rect 12378 19276 12394 19444
rect 12428 19276 12466 19444
rect 12378 19260 12466 19276
rect 13266 19444 13354 19460
rect 13266 19276 13304 19444
rect 13338 19276 13354 19444
rect 13266 19260 13354 19276
rect 13859 19444 13947 19460
rect 13859 19276 13875 19444
rect 13909 19276 13947 19444
rect 13859 19260 13947 19276
rect 14747 19444 14835 19460
rect 14747 19276 14785 19444
rect 14819 19276 14835 19444
rect 14747 19260 14835 19276
rect 12378 19186 12466 19202
rect 12378 19018 12394 19186
rect 12428 19018 12466 19186
rect 12378 19002 12466 19018
rect 13266 19186 13354 19202
rect 13266 19018 13304 19186
rect 13338 19018 13354 19186
rect 13266 19002 13354 19018
rect 13859 19186 13947 19202
rect 13859 19018 13875 19186
rect 13909 19018 13947 19186
rect 13859 19002 13947 19018
rect 14747 19186 14835 19202
rect 14747 19018 14785 19186
rect 14819 19018 14835 19186
rect 14747 19002 14835 19018
rect 12378 18928 12466 18944
rect 12378 18760 12394 18928
rect 12428 18760 12466 18928
rect 12378 18744 12466 18760
rect 13266 18928 13354 18944
rect 13266 18760 13304 18928
rect 13338 18760 13354 18928
rect 13266 18744 13354 18760
rect 13859 18928 13947 18944
rect 13859 18760 13875 18928
rect 13909 18760 13947 18928
rect 13859 18744 13947 18760
rect 14747 18928 14835 18944
rect 14747 18760 14785 18928
rect 14819 18760 14835 18928
rect 14747 18744 14835 18760
rect 12378 18670 12466 18686
rect 12378 18502 12394 18670
rect 12428 18502 12466 18670
rect 12378 18486 12466 18502
rect 13266 18670 13354 18686
rect 13266 18502 13304 18670
rect 13338 18502 13354 18670
rect 13266 18486 13354 18502
rect 13859 18670 13947 18686
rect 13859 18502 13875 18670
rect 13909 18502 13947 18670
rect 13859 18486 13947 18502
rect 14747 18670 14835 18686
rect 14747 18502 14785 18670
rect 14819 18502 14835 18670
rect 14747 18486 14835 18502
rect 12378 18412 12466 18428
rect 12378 18244 12394 18412
rect 12428 18244 12466 18412
rect 12378 18228 12466 18244
rect 13266 18412 13354 18428
rect 13266 18244 13304 18412
rect 13338 18244 13354 18412
rect 13266 18228 13354 18244
rect 13859 18412 13947 18428
rect 13859 18244 13875 18412
rect 13909 18244 13947 18412
rect 13859 18228 13947 18244
rect 14747 18412 14835 18428
rect 14747 18244 14785 18412
rect 14819 18244 14835 18412
rect 14747 18228 14835 18244
rect 12378 18154 12466 18170
rect 12378 17986 12394 18154
rect 12428 17986 12466 18154
rect 12378 17970 12466 17986
rect 13266 18154 13354 18170
rect 13266 17986 13304 18154
rect 13338 17986 13354 18154
rect 13266 17970 13354 17986
rect 13859 18154 13947 18170
rect 13859 17986 13875 18154
rect 13909 17986 13947 18154
rect 13859 17970 13947 17986
rect 14747 18154 14835 18170
rect 14747 17986 14785 18154
rect 14819 17986 14835 18154
rect 14747 17970 14835 17986
rect 12378 17896 12466 17912
rect 12378 17728 12394 17896
rect 12428 17728 12466 17896
rect 12378 17712 12466 17728
rect 13266 17896 13354 17912
rect 13266 17728 13304 17896
rect 13338 17728 13354 17896
rect 13266 17712 13354 17728
rect 13859 17896 13947 17912
rect 13859 17728 13875 17896
rect 13909 17728 13947 17896
rect 13859 17712 13947 17728
rect 14747 17896 14835 17912
rect 14747 17728 14785 17896
rect 14819 17728 14835 17896
rect 14747 17712 14835 17728
rect 12378 17638 12466 17654
rect 12378 17470 12394 17638
rect 12428 17470 12466 17638
rect 12378 17454 12466 17470
rect 13266 17638 13354 17654
rect 13266 17470 13304 17638
rect 13338 17470 13354 17638
rect 13266 17454 13354 17470
rect 13859 17638 13947 17654
rect 13859 17470 13875 17638
rect 13909 17470 13947 17638
rect 13859 17454 13947 17470
rect 14747 17638 14835 17654
rect 14747 17470 14785 17638
rect 14819 17470 14835 17638
rect 14747 17454 14835 17470
rect 12378 17380 12466 17396
rect 12378 17212 12394 17380
rect 12428 17212 12466 17380
rect 12378 17196 12466 17212
rect 13266 17380 13354 17396
rect 13266 17212 13304 17380
rect 13338 17212 13354 17380
rect 13266 17196 13354 17212
rect 13859 17380 13947 17396
rect 13859 17212 13875 17380
rect 13909 17212 13947 17380
rect 13859 17196 13947 17212
rect 14747 17380 14835 17396
rect 14747 17212 14785 17380
rect 14819 17212 14835 17380
rect 14747 17196 14835 17212
rect 12378 17122 12466 17138
rect 12378 16954 12394 17122
rect 12428 16954 12466 17122
rect 12378 16938 12466 16954
rect 13266 17122 13354 17138
rect 13266 16954 13304 17122
rect 13338 16954 13354 17122
rect 13266 16938 13354 16954
rect 13859 17122 13947 17138
rect 13859 16954 13875 17122
rect 13909 16954 13947 17122
rect 13859 16938 13947 16954
rect 14747 17122 14835 17138
rect 14747 16954 14785 17122
rect 14819 16954 14835 17122
rect 14747 16938 14835 16954
rect 12378 16864 12466 16880
rect 12378 16696 12394 16864
rect 12428 16696 12466 16864
rect 12378 16680 12466 16696
rect 13266 16864 13354 16880
rect 13266 16696 13304 16864
rect 13338 16696 13354 16864
rect 13266 16680 13354 16696
rect 13859 16864 13947 16880
rect 13859 16696 13875 16864
rect 13909 16696 13947 16864
rect 13859 16680 13947 16696
rect 14747 16864 14835 16880
rect 14747 16696 14785 16864
rect 14819 16696 14835 16864
rect 14747 16680 14835 16696
rect 12378 16606 12466 16622
rect 12378 16438 12394 16606
rect 12428 16438 12466 16606
rect 12378 16422 12466 16438
rect 13266 16606 13354 16622
rect 13266 16438 13304 16606
rect 13338 16438 13354 16606
rect 13266 16422 13354 16438
rect 13859 16606 13947 16622
rect 13859 16438 13875 16606
rect 13909 16438 13947 16606
rect 13859 16422 13947 16438
rect 14747 16606 14835 16622
rect 14747 16438 14785 16606
rect 14819 16438 14835 16606
rect 14747 16422 14835 16438
rect 12378 16348 12466 16364
rect 12378 16180 12394 16348
rect 12428 16180 12466 16348
rect 12378 16164 12466 16180
rect 13266 16348 13354 16364
rect 13266 16180 13304 16348
rect 13338 16180 13354 16348
rect 13266 16164 13354 16180
rect 13859 16348 13947 16364
rect 13859 16180 13875 16348
rect 13909 16180 13947 16348
rect 13859 16164 13947 16180
rect 14747 16348 14835 16364
rect 14747 16180 14785 16348
rect 14819 16180 14835 16348
rect 14747 16164 14835 16180
rect 12378 16090 12466 16106
rect 12378 15922 12394 16090
rect 12428 15922 12466 16090
rect 12378 15906 12466 15922
rect 13266 16090 13354 16106
rect 13266 15922 13304 16090
rect 13338 15922 13354 16090
rect 13266 15906 13354 15922
rect 13859 16090 13947 16106
rect 13859 15922 13875 16090
rect 13909 15922 13947 16090
rect 13859 15906 13947 15922
rect 14747 16090 14835 16106
rect 14747 15922 14785 16090
rect 14819 15922 14835 16090
rect 14747 15906 14835 15922
rect 12378 15832 12466 15848
rect 12378 15664 12394 15832
rect 12428 15664 12466 15832
rect 12378 15648 12466 15664
rect 13266 15832 13354 15848
rect 13266 15664 13304 15832
rect 13338 15664 13354 15832
rect 13266 15648 13354 15664
rect 13859 15832 13947 15848
rect 13859 15664 13875 15832
rect 13909 15664 13947 15832
rect 13859 15648 13947 15664
rect 14747 15832 14835 15848
rect 14747 15664 14785 15832
rect 14819 15664 14835 15832
rect 14747 15648 14835 15664
rect 12378 15574 12466 15590
rect 12378 15406 12394 15574
rect 12428 15406 12466 15574
rect 12378 15390 12466 15406
rect 13266 15574 13354 15590
rect 13266 15406 13304 15574
rect 13338 15406 13354 15574
rect 13266 15390 13354 15406
rect 13859 15574 13947 15590
rect 13859 15406 13875 15574
rect 13909 15406 13947 15574
rect 13859 15390 13947 15406
rect 14747 15574 14835 15590
rect 14747 15406 14785 15574
rect 14819 15406 14835 15574
rect 14747 15390 14835 15406
rect 15996 22313 16084 22329
rect 15996 22145 16012 22313
rect 16046 22145 16084 22313
rect 15996 22129 16084 22145
rect 16284 22313 16372 22329
rect 16284 22145 16322 22313
rect 16356 22145 16372 22313
rect 16284 22129 16372 22145
rect 15996 22055 16084 22071
rect 15996 21887 16012 22055
rect 16046 21887 16084 22055
rect 15996 21871 16084 21887
rect 16284 22055 16372 22071
rect 16284 21887 16322 22055
rect 16356 21887 16372 22055
rect 16284 21871 16372 21887
rect 15996 21797 16084 21813
rect 15996 21629 16012 21797
rect 16046 21629 16084 21797
rect 15996 21613 16084 21629
rect 16284 21797 16372 21813
rect 16284 21629 16322 21797
rect 16356 21629 16372 21797
rect 16284 21613 16372 21629
rect 15996 21539 16084 21555
rect 15996 21371 16012 21539
rect 16046 21371 16084 21539
rect 15996 21355 16084 21371
rect 16284 21539 16372 21555
rect 16284 21371 16322 21539
rect 16356 21371 16372 21539
rect 16284 21355 16372 21371
rect 15996 21281 16084 21297
rect 15996 21113 16012 21281
rect 16046 21113 16084 21281
rect 15996 21097 16084 21113
rect 16284 21281 16372 21297
rect 16284 21113 16322 21281
rect 16356 21113 16372 21281
rect 16284 21097 16372 21113
rect 15996 21023 16084 21039
rect 15996 20855 16012 21023
rect 16046 20855 16084 21023
rect 15996 20839 16084 20855
rect 16284 21023 16372 21039
rect 16284 20855 16322 21023
rect 16356 20855 16372 21023
rect 16284 20839 16372 20855
rect 15996 20765 16084 20781
rect 15996 20597 16012 20765
rect 16046 20597 16084 20765
rect 15996 20581 16084 20597
rect 16284 20765 16372 20781
rect 16284 20597 16322 20765
rect 16356 20597 16372 20765
rect 16284 20581 16372 20597
rect 15996 20507 16084 20523
rect 15996 20339 16012 20507
rect 16046 20339 16084 20507
rect 15996 20323 16084 20339
rect 16284 20507 16372 20523
rect 16284 20339 16322 20507
rect 16356 20339 16372 20507
rect 16284 20323 16372 20339
rect 15996 20249 16084 20265
rect 15996 20081 16012 20249
rect 16046 20081 16084 20249
rect 15996 20065 16084 20081
rect 16284 20249 16372 20265
rect 16284 20081 16322 20249
rect 16356 20081 16372 20249
rect 16284 20065 16372 20081
rect 15996 19991 16084 20007
rect 15996 19823 16012 19991
rect 16046 19823 16084 19991
rect 15996 19807 16084 19823
rect 16284 19991 16372 20007
rect 16284 19823 16322 19991
rect 16356 19823 16372 19991
rect 16284 19807 16372 19823
rect 15996 19733 16084 19749
rect 15996 19565 16012 19733
rect 16046 19565 16084 19733
rect 15996 19549 16084 19565
rect 16284 19733 16372 19749
rect 16284 19565 16322 19733
rect 16356 19565 16372 19733
rect 16284 19549 16372 19565
rect 15996 19475 16084 19491
rect 15996 19307 16012 19475
rect 16046 19307 16084 19475
rect 15996 19291 16084 19307
rect 16284 19475 16372 19491
rect 16284 19307 16322 19475
rect 16356 19307 16372 19475
rect 16284 19291 16372 19307
rect 15996 19217 16084 19233
rect 15996 19049 16012 19217
rect 16046 19049 16084 19217
rect 15996 19033 16084 19049
rect 16284 19217 16372 19233
rect 16284 19049 16322 19217
rect 16356 19049 16372 19217
rect 16284 19033 16372 19049
rect 15996 18959 16084 18975
rect 15996 18791 16012 18959
rect 16046 18791 16084 18959
rect 15996 18775 16084 18791
rect 16284 18959 16372 18975
rect 16284 18791 16322 18959
rect 16356 18791 16372 18959
rect 16284 18775 16372 18791
rect 15996 18701 16084 18717
rect 15996 18533 16012 18701
rect 16046 18533 16084 18701
rect 15996 18517 16084 18533
rect 16284 18701 16372 18717
rect 16284 18533 16322 18701
rect 16356 18533 16372 18701
rect 16284 18517 16372 18533
rect 15996 18443 16084 18459
rect 15996 18275 16012 18443
rect 16046 18275 16084 18443
rect 15996 18259 16084 18275
rect 16284 18443 16372 18459
rect 16284 18275 16322 18443
rect 16356 18275 16372 18443
rect 16284 18259 16372 18275
rect 15996 18185 16084 18201
rect 15996 18017 16012 18185
rect 16046 18017 16084 18185
rect 15996 18001 16084 18017
rect 16284 18185 16372 18201
rect 16284 18017 16322 18185
rect 16356 18017 16372 18185
rect 16284 18001 16372 18017
rect 15996 17927 16084 17943
rect 15996 17759 16012 17927
rect 16046 17759 16084 17927
rect 15996 17743 16084 17759
rect 16284 17927 16372 17943
rect 16284 17759 16322 17927
rect 16356 17759 16372 17927
rect 16284 17743 16372 17759
rect 15996 17669 16084 17685
rect 15996 17501 16012 17669
rect 16046 17501 16084 17669
rect 15996 17485 16084 17501
rect 16284 17669 16372 17685
rect 16284 17501 16322 17669
rect 16356 17501 16372 17669
rect 16284 17485 16372 17501
rect 15996 17411 16084 17427
rect 15996 17243 16012 17411
rect 16046 17243 16084 17411
rect 15996 17227 16084 17243
rect 16284 17411 16372 17427
rect 16284 17243 16322 17411
rect 16356 17243 16372 17411
rect 16284 17227 16372 17243
rect 16774 22378 16871 22394
rect 16774 22010 16790 22378
rect 16824 22010 16871 22378
rect 16774 21994 16871 22010
rect 17071 22378 17168 22394
rect 17071 22010 17118 22378
rect 17152 22010 17168 22378
rect 17071 21994 17168 22010
rect 16774 21797 16871 21813
rect 16774 21429 16790 21797
rect 16824 21429 16871 21797
rect 16774 21413 16871 21429
rect 17071 21797 17168 21813
rect 17071 21429 17118 21797
rect 17152 21429 17168 21797
rect 17071 21413 17168 21429
rect 22566 22688 22654 22704
rect 22566 22420 22582 22688
rect 22616 22420 22654 22688
rect 22566 22404 22654 22420
rect 23754 22688 23842 22704
rect 23754 22420 23792 22688
rect 23826 22420 23842 22688
rect 23754 22404 23842 22420
rect 22566 22330 22654 22346
rect 22566 22062 22582 22330
rect 22616 22062 22654 22330
rect 22566 22046 22654 22062
rect 23754 22330 23842 22346
rect 23754 22062 23792 22330
rect 23826 22062 23842 22330
rect 23754 22046 23842 22062
rect 16774 20507 16871 20523
rect 16774 20139 16790 20507
rect 16824 20139 16871 20507
rect 16774 20123 16871 20139
rect 17071 20507 17168 20523
rect 17071 20139 17118 20507
rect 17152 20139 17168 20507
rect 17071 20123 17168 20139
rect 16774 19217 16871 19233
rect 16774 18849 16790 19217
rect 16824 18849 16871 19217
rect 16774 18833 16871 18849
rect 17071 19217 17168 19233
rect 17071 18849 17118 19217
rect 17152 18849 17168 19217
rect 17071 18833 17168 18849
rect 16774 17927 16871 17943
rect 16774 17559 16790 17927
rect 16824 17559 16871 17927
rect 16774 17543 16871 17559
rect 17071 17927 17168 17943
rect 17071 17559 17118 17927
rect 17152 17559 17168 17927
rect 17071 17543 17168 17559
rect 16774 16839 16871 16855
rect 16774 16671 16790 16839
rect 16824 16671 16871 16839
rect 16774 16655 16871 16671
rect 17071 16839 17168 16855
rect 17071 16671 17118 16839
rect 17152 16671 17168 16839
rect 17071 16655 17168 16671
rect 16774 16581 16871 16597
rect 16774 16413 16790 16581
rect 16824 16413 16871 16581
rect 16774 16397 16871 16413
rect 17071 16581 17168 16597
rect 17071 16413 17118 16581
rect 17152 16413 17168 16581
rect 17071 16397 17168 16413
rect 16774 16114 16871 16130
rect 16774 15746 16790 16114
rect 16824 15746 16871 16114
rect 16774 15730 16871 15746
rect 16971 16114 17068 16130
rect 16971 15746 17018 16114
rect 17052 15746 17068 16114
rect 16971 15730 17068 15746
rect 16774 15656 16871 15672
rect 16774 15288 16790 15656
rect 16824 15288 16871 15656
rect 16774 15272 16871 15288
rect 16971 15656 17068 15672
rect 16971 15288 17018 15656
rect 17052 15288 17068 15656
rect 16971 15272 17068 15288
rect 3013 10123 3101 10139
rect 3013 9955 3029 10123
rect 3063 9955 3101 10123
rect 3013 9939 3101 9955
rect 3901 10123 3989 10139
rect 3901 9955 3939 10123
rect 3973 9955 3989 10123
rect 3901 9939 3989 9955
rect 4494 10123 4582 10139
rect 4494 9955 4510 10123
rect 4544 9955 4582 10123
rect 4494 9939 4582 9955
rect 5382 10123 5470 10139
rect 5382 9955 5420 10123
rect 5454 9955 5470 10123
rect 5382 9939 5470 9955
rect 3013 9865 3101 9881
rect 3013 9697 3029 9865
rect 3063 9697 3101 9865
rect 3013 9681 3101 9697
rect 3901 9865 3989 9881
rect 3901 9697 3939 9865
rect 3973 9697 3989 9865
rect 3901 9681 3989 9697
rect 4494 9865 4582 9881
rect 4494 9697 4510 9865
rect 4544 9697 4582 9865
rect 4494 9681 4582 9697
rect 5382 9865 5470 9881
rect 5382 9697 5420 9865
rect 5454 9697 5470 9865
rect 5382 9681 5470 9697
rect 3013 9607 3101 9623
rect 3013 9439 3029 9607
rect 3063 9439 3101 9607
rect 3013 9423 3101 9439
rect 3901 9607 3989 9623
rect 3901 9439 3939 9607
rect 3973 9439 3989 9607
rect 3901 9423 3989 9439
rect 4494 9607 4582 9623
rect 4494 9439 4510 9607
rect 4544 9439 4582 9607
rect 4494 9423 4582 9439
rect 5382 9607 5470 9623
rect 5382 9439 5420 9607
rect 5454 9439 5470 9607
rect 5382 9423 5470 9439
rect 3013 9349 3101 9365
rect 3013 9181 3029 9349
rect 3063 9181 3101 9349
rect 3013 9165 3101 9181
rect 3901 9349 3989 9365
rect 3901 9181 3939 9349
rect 3973 9181 3989 9349
rect 3901 9165 3989 9181
rect 4494 9349 4582 9365
rect 4494 9181 4510 9349
rect 4544 9181 4582 9349
rect 4494 9165 4582 9181
rect 5382 9349 5470 9365
rect 5382 9181 5420 9349
rect 5454 9181 5470 9349
rect 5382 9165 5470 9181
rect 3013 9091 3101 9107
rect 3013 8923 3029 9091
rect 3063 8923 3101 9091
rect 3013 8907 3101 8923
rect 3901 9091 3989 9107
rect 3901 8923 3939 9091
rect 3973 8923 3989 9091
rect 3901 8907 3989 8923
rect 4494 9091 4582 9107
rect 4494 8923 4510 9091
rect 4544 8923 4582 9091
rect 4494 8907 4582 8923
rect 5382 9091 5470 9107
rect 5382 8923 5420 9091
rect 5454 8923 5470 9091
rect 5382 8907 5470 8923
rect 3013 8833 3101 8849
rect 3013 8665 3029 8833
rect 3063 8665 3101 8833
rect 3013 8649 3101 8665
rect 3901 8833 3989 8849
rect 3901 8665 3939 8833
rect 3973 8665 3989 8833
rect 3901 8649 3989 8665
rect 4494 8833 4582 8849
rect 4494 8665 4510 8833
rect 4544 8665 4582 8833
rect 4494 8649 4582 8665
rect 5382 8833 5470 8849
rect 5382 8665 5420 8833
rect 5454 8665 5470 8833
rect 5382 8649 5470 8665
rect 3013 8575 3101 8591
rect 3013 8407 3029 8575
rect 3063 8407 3101 8575
rect 3013 8391 3101 8407
rect 3901 8575 3989 8591
rect 3901 8407 3939 8575
rect 3973 8407 3989 8575
rect 3901 8391 3989 8407
rect 4494 8575 4582 8591
rect 4494 8407 4510 8575
rect 4544 8407 4582 8575
rect 4494 8391 4582 8407
rect 5382 8575 5470 8591
rect 5382 8407 5420 8575
rect 5454 8407 5470 8575
rect 5382 8391 5470 8407
rect 3013 8317 3101 8333
rect 3013 8149 3029 8317
rect 3063 8149 3101 8317
rect 3013 8133 3101 8149
rect 3901 8317 3989 8333
rect 3901 8149 3939 8317
rect 3973 8149 3989 8317
rect 3901 8133 3989 8149
rect 4494 8317 4582 8333
rect 4494 8149 4510 8317
rect 4544 8149 4582 8317
rect 4494 8133 4582 8149
rect 5382 8317 5470 8333
rect 5382 8149 5420 8317
rect 5454 8149 5470 8317
rect 5382 8133 5470 8149
rect 3013 8059 3101 8075
rect 3013 7891 3029 8059
rect 3063 7891 3101 8059
rect 3013 7875 3101 7891
rect 3901 8059 3989 8075
rect 3901 7891 3939 8059
rect 3973 7891 3989 8059
rect 3901 7875 3989 7891
rect 4494 8059 4582 8075
rect 4494 7891 4510 8059
rect 4544 7891 4582 8059
rect 4494 7875 4582 7891
rect 5382 8059 5470 8075
rect 5382 7891 5420 8059
rect 5454 7891 5470 8059
rect 5382 7875 5470 7891
rect 3013 7801 3101 7817
rect 3013 7633 3029 7801
rect 3063 7633 3101 7801
rect 3013 7617 3101 7633
rect 3901 7801 3989 7817
rect 3901 7633 3939 7801
rect 3973 7633 3989 7801
rect 3901 7617 3989 7633
rect 4494 7801 4582 7817
rect 4494 7633 4510 7801
rect 4544 7633 4582 7801
rect 4494 7617 4582 7633
rect 5382 7801 5470 7817
rect 5382 7633 5420 7801
rect 5454 7633 5470 7801
rect 5382 7617 5470 7633
rect 3013 7543 3101 7559
rect 3013 7375 3029 7543
rect 3063 7375 3101 7543
rect 3013 7359 3101 7375
rect 3901 7543 3989 7559
rect 3901 7375 3939 7543
rect 3973 7375 3989 7543
rect 3901 7359 3989 7375
rect 4494 7543 4582 7559
rect 4494 7375 4510 7543
rect 4544 7375 4582 7543
rect 4494 7359 4582 7375
rect 5382 7543 5470 7559
rect 5382 7375 5420 7543
rect 5454 7375 5470 7543
rect 5382 7359 5470 7375
rect 3013 7285 3101 7301
rect 3013 7117 3029 7285
rect 3063 7117 3101 7285
rect 3013 7101 3101 7117
rect 3901 7285 3989 7301
rect 3901 7117 3939 7285
rect 3973 7117 3989 7285
rect 3901 7101 3989 7117
rect 4494 7285 4582 7301
rect 4494 7117 4510 7285
rect 4544 7117 4582 7285
rect 4494 7101 4582 7117
rect 5382 7285 5470 7301
rect 5382 7117 5420 7285
rect 5454 7117 5470 7285
rect 5382 7101 5470 7117
rect 3013 7027 3101 7043
rect 3013 6859 3029 7027
rect 3063 6859 3101 7027
rect 3013 6843 3101 6859
rect 3901 7027 3989 7043
rect 3901 6859 3939 7027
rect 3973 6859 3989 7027
rect 3901 6843 3989 6859
rect 4494 7027 4582 7043
rect 4494 6859 4510 7027
rect 4544 6859 4582 7027
rect 4494 6843 4582 6859
rect 5382 7027 5470 7043
rect 5382 6859 5420 7027
rect 5454 6859 5470 7027
rect 5382 6843 5470 6859
rect 3013 6769 3101 6785
rect 3013 6601 3029 6769
rect 3063 6601 3101 6769
rect 3013 6585 3101 6601
rect 3901 6769 3989 6785
rect 3901 6601 3939 6769
rect 3973 6601 3989 6769
rect 3901 6585 3989 6601
rect 4494 6769 4582 6785
rect 4494 6601 4510 6769
rect 4544 6601 4582 6769
rect 4494 6585 4582 6601
rect 5382 6769 5470 6785
rect 5382 6601 5420 6769
rect 5454 6601 5470 6769
rect 5382 6585 5470 6601
rect 3013 6511 3101 6527
rect 3013 6343 3029 6511
rect 3063 6343 3101 6511
rect 3013 6327 3101 6343
rect 3901 6511 3989 6527
rect 3901 6343 3939 6511
rect 3973 6343 3989 6511
rect 3901 6327 3989 6343
rect 4494 6511 4582 6527
rect 4494 6343 4510 6511
rect 4544 6343 4582 6511
rect 4494 6327 4582 6343
rect 5382 6511 5470 6527
rect 5382 6343 5420 6511
rect 5454 6343 5470 6511
rect 5382 6327 5470 6343
rect 3013 6253 3101 6269
rect 3013 6085 3029 6253
rect 3063 6085 3101 6253
rect 3013 6069 3101 6085
rect 3901 6253 3989 6269
rect 3901 6085 3939 6253
rect 3973 6085 3989 6253
rect 3901 6069 3989 6085
rect 4494 6253 4582 6269
rect 4494 6085 4510 6253
rect 4544 6085 4582 6253
rect 4494 6069 4582 6085
rect 5382 6253 5470 6269
rect 5382 6085 5420 6253
rect 5454 6085 5470 6253
rect 5382 6069 5470 6085
rect 3013 5995 3101 6011
rect 3013 5827 3029 5995
rect 3063 5827 3101 5995
rect 3013 5811 3101 5827
rect 3901 5995 3989 6011
rect 3901 5827 3939 5995
rect 3973 5827 3989 5995
rect 3901 5811 3989 5827
rect 4494 5995 4582 6011
rect 4494 5827 4510 5995
rect 4544 5827 4582 5995
rect 4494 5811 4582 5827
rect 5382 5995 5470 6011
rect 5382 5827 5420 5995
rect 5454 5827 5470 5995
rect 5382 5811 5470 5827
rect 3013 5737 3101 5753
rect 3013 5569 3029 5737
rect 3063 5569 3101 5737
rect 3013 5553 3101 5569
rect 3901 5737 3989 5753
rect 3901 5569 3939 5737
rect 3973 5569 3989 5737
rect 3901 5553 3989 5569
rect 4494 5737 4582 5753
rect 4494 5569 4510 5737
rect 4544 5569 4582 5737
rect 4494 5553 4582 5569
rect 5382 5737 5470 5753
rect 5382 5569 5420 5737
rect 5454 5569 5470 5737
rect 5382 5553 5470 5569
rect 3013 5479 3101 5495
rect 3013 5311 3029 5479
rect 3063 5311 3101 5479
rect 3013 5295 3101 5311
rect 3901 5479 3989 5495
rect 3901 5311 3939 5479
rect 3973 5311 3989 5479
rect 3901 5295 3989 5311
rect 4494 5479 4582 5495
rect 4494 5311 4510 5479
rect 4544 5311 4582 5479
rect 4494 5295 4582 5311
rect 5382 5479 5470 5495
rect 5382 5311 5420 5479
rect 5454 5311 5470 5479
rect 5382 5295 5470 5311
rect 3013 5221 3101 5237
rect 3013 5053 3029 5221
rect 3063 5053 3101 5221
rect 3013 5037 3101 5053
rect 3901 5221 3989 5237
rect 3901 5053 3939 5221
rect 3973 5053 3989 5221
rect 3901 5037 3989 5053
rect 4494 5221 4582 5237
rect 4494 5053 4510 5221
rect 4544 5053 4582 5221
rect 4494 5037 4582 5053
rect 5382 5221 5470 5237
rect 5382 5053 5420 5221
rect 5454 5053 5470 5221
rect 5382 5037 5470 5053
rect 3013 4963 3101 4979
rect 3013 4795 3029 4963
rect 3063 4795 3101 4963
rect 3013 4779 3101 4795
rect 3901 4963 3989 4979
rect 3901 4795 3939 4963
rect 3973 4795 3989 4963
rect 3901 4779 3989 4795
rect 4494 4963 4582 4979
rect 4494 4795 4510 4963
rect 4544 4795 4582 4963
rect 4494 4779 4582 4795
rect 5382 4963 5470 4979
rect 5382 4795 5420 4963
rect 5454 4795 5470 4963
rect 5382 4779 5470 4795
rect 3013 4705 3101 4721
rect 3013 4537 3029 4705
rect 3063 4537 3101 4705
rect 3013 4521 3101 4537
rect 3901 4705 3989 4721
rect 3901 4537 3939 4705
rect 3973 4537 3989 4705
rect 3901 4521 3989 4537
rect 4494 4705 4582 4721
rect 4494 4537 4510 4705
rect 4544 4537 4582 4705
rect 4494 4521 4582 4537
rect 5382 4705 5470 4721
rect 5382 4537 5420 4705
rect 5454 4537 5470 4705
rect 5382 4521 5470 4537
rect 3013 4447 3101 4463
rect 3013 4279 3029 4447
rect 3063 4279 3101 4447
rect 3013 4263 3101 4279
rect 3901 4447 3989 4463
rect 3901 4279 3939 4447
rect 3973 4279 3989 4447
rect 3901 4263 3989 4279
rect 4494 4447 4582 4463
rect 4494 4279 4510 4447
rect 4544 4279 4582 4447
rect 4494 4263 4582 4279
rect 5382 4447 5470 4463
rect 5382 4279 5420 4447
rect 5454 4279 5470 4447
rect 5382 4263 5470 4279
rect 3013 4189 3101 4205
rect 3013 4021 3029 4189
rect 3063 4021 3101 4189
rect 3013 4005 3101 4021
rect 3901 4189 3989 4205
rect 3901 4021 3939 4189
rect 3973 4021 3989 4189
rect 3901 4005 3989 4021
rect 4494 4189 4582 4205
rect 4494 4021 4510 4189
rect 4544 4021 4582 4189
rect 4494 4005 4582 4021
rect 5382 4189 5470 4205
rect 5382 4021 5420 4189
rect 5454 4021 5470 4189
rect 5382 4005 5470 4021
rect 7409 10241 7506 10257
rect 7409 9873 7425 10241
rect 7459 9873 7506 10241
rect 7409 9857 7506 9873
rect 7606 10241 7703 10257
rect 7606 9873 7653 10241
rect 7687 9873 7703 10241
rect 7606 9857 7703 9873
rect 7409 9783 7506 9799
rect 7409 9415 7425 9783
rect 7459 9415 7506 9783
rect 7409 9399 7506 9415
rect 7606 9783 7703 9799
rect 7606 9415 7653 9783
rect 7687 9415 7703 9783
rect 7606 9399 7703 9415
rect 7409 9116 7506 9132
rect 7409 8948 7425 9116
rect 7459 8948 7506 9116
rect 7409 8932 7506 8948
rect 7706 9116 7803 9132
rect 7706 8948 7753 9116
rect 7787 8948 7803 9116
rect 7706 8932 7803 8948
rect 7409 8858 7506 8874
rect 7409 8690 7425 8858
rect 7459 8690 7506 8858
rect 7409 8674 7506 8690
rect 7706 8858 7803 8874
rect 7706 8690 7753 8858
rect 7787 8690 7803 8858
rect 7706 8674 7803 8690
rect 18221 10747 21821 10763
rect 18221 10713 18237 10747
rect 21805 10713 21821 10747
rect 18221 10666 21821 10713
rect 21879 10747 25479 10763
rect 21879 10713 21895 10747
rect 25463 10713 25479 10747
rect 21879 10666 25479 10713
rect 18221 10259 21821 10306
rect 18221 10225 18237 10259
rect 21805 10225 21821 10259
rect 18221 10178 21821 10225
rect 21879 10259 25479 10306
rect 21879 10225 21895 10259
rect 25463 10225 25479 10259
rect 21879 10178 25479 10225
rect 18221 9771 21821 9818
rect 18221 9737 18237 9771
rect 21805 9737 21821 9771
rect 18221 9721 21821 9737
rect 21879 9771 25479 9818
rect 21879 9737 21895 9771
rect 25463 9737 25479 9771
rect 21879 9721 25479 9737
rect 6631 8187 6719 8203
rect 6631 8019 6647 8187
rect 6681 8019 6719 8187
rect 6631 8003 6719 8019
rect 6919 8187 7007 8203
rect 6919 8019 6957 8187
rect 6991 8019 7007 8187
rect 6919 8003 7007 8019
rect 6631 7929 6719 7945
rect 6631 7761 6647 7929
rect 6681 7761 6719 7929
rect 6631 7745 6719 7761
rect 6919 7929 7007 7945
rect 6919 7761 6957 7929
rect 6991 7761 7007 7929
rect 6919 7745 7007 7761
rect 6631 7671 6719 7687
rect 6631 7503 6647 7671
rect 6681 7503 6719 7671
rect 6631 7487 6719 7503
rect 6919 7671 7007 7687
rect 6919 7503 6957 7671
rect 6991 7503 7007 7671
rect 6919 7487 7007 7503
rect 6631 7413 6719 7429
rect 6631 7245 6647 7413
rect 6681 7245 6719 7413
rect 6631 7229 6719 7245
rect 6919 7413 7007 7429
rect 6919 7245 6957 7413
rect 6991 7245 7007 7413
rect 6919 7229 7007 7245
rect 6631 7155 6719 7171
rect 6631 6987 6647 7155
rect 6681 6987 6719 7155
rect 6631 6971 6719 6987
rect 6919 7155 7007 7171
rect 6919 6987 6957 7155
rect 6991 6987 7007 7155
rect 6919 6971 7007 6987
rect 6631 6897 6719 6913
rect 6631 6729 6647 6897
rect 6681 6729 6719 6897
rect 6631 6713 6719 6729
rect 6919 6897 7007 6913
rect 6919 6729 6957 6897
rect 6991 6729 7007 6897
rect 6919 6713 7007 6729
rect 6631 6639 6719 6655
rect 6631 6471 6647 6639
rect 6681 6471 6719 6639
rect 6631 6455 6719 6471
rect 6919 6639 7007 6655
rect 6919 6471 6957 6639
rect 6991 6471 7007 6639
rect 6919 6455 7007 6471
rect 6631 6381 6719 6397
rect 6631 6213 6647 6381
rect 6681 6213 6719 6381
rect 6631 6197 6719 6213
rect 6919 6381 7007 6397
rect 6919 6213 6957 6381
rect 6991 6213 7007 6381
rect 6919 6197 7007 6213
rect 6631 6123 6719 6139
rect 6631 5955 6647 6123
rect 6681 5955 6719 6123
rect 6631 5939 6719 5955
rect 6919 6123 7007 6139
rect 6919 5955 6957 6123
rect 6991 5955 7007 6123
rect 6919 5939 7007 5955
rect 6631 5865 6719 5881
rect 6631 5697 6647 5865
rect 6681 5697 6719 5865
rect 6631 5681 6719 5697
rect 6919 5865 7007 5881
rect 6919 5697 6957 5865
rect 6991 5697 7007 5865
rect 6919 5681 7007 5697
rect 6631 5607 6719 5623
rect 6631 5439 6647 5607
rect 6681 5439 6719 5607
rect 6631 5423 6719 5439
rect 6919 5607 7007 5623
rect 6919 5439 6957 5607
rect 6991 5439 7007 5607
rect 6919 5423 7007 5439
rect 6631 5349 6719 5365
rect 6631 5181 6647 5349
rect 6681 5181 6719 5349
rect 6631 5165 6719 5181
rect 6919 5349 7007 5365
rect 6919 5181 6957 5349
rect 6991 5181 7007 5349
rect 6919 5165 7007 5181
rect 6631 5091 6719 5107
rect 6631 4923 6647 5091
rect 6681 4923 6719 5091
rect 6631 4907 6719 4923
rect 6919 5091 7007 5107
rect 6919 4923 6957 5091
rect 6991 4923 7007 5091
rect 6919 4907 7007 4923
rect 6631 4833 6719 4849
rect 6631 4665 6647 4833
rect 6681 4665 6719 4833
rect 6631 4649 6719 4665
rect 6919 4833 7007 4849
rect 6919 4665 6957 4833
rect 6991 4665 7007 4833
rect 6919 4649 7007 4665
rect 6631 4575 6719 4591
rect 6631 4407 6647 4575
rect 6681 4407 6719 4575
rect 6631 4391 6719 4407
rect 6919 4575 7007 4591
rect 6919 4407 6957 4575
rect 6991 4407 7007 4575
rect 6919 4391 7007 4407
rect 6631 4317 6719 4333
rect 6631 4149 6647 4317
rect 6681 4149 6719 4317
rect 6631 4133 6719 4149
rect 6919 4317 7007 4333
rect 6919 4149 6957 4317
rect 6991 4149 7007 4317
rect 6919 4133 7007 4149
rect 6631 4059 6719 4075
rect 6631 3891 6647 4059
rect 6681 3891 6719 4059
rect 6631 3875 6719 3891
rect 6919 4059 7007 4075
rect 6919 3891 6957 4059
rect 6991 3891 7007 4059
rect 6919 3875 7007 3891
rect 6631 3801 6719 3817
rect 6631 3633 6647 3801
rect 6681 3633 6719 3801
rect 6631 3617 6719 3633
rect 6919 3801 7007 3817
rect 6919 3633 6957 3801
rect 6991 3633 7007 3801
rect 6919 3617 7007 3633
rect 6631 3543 6719 3559
rect 6631 3375 6647 3543
rect 6681 3375 6719 3543
rect 6631 3359 6719 3375
rect 6919 3543 7007 3559
rect 6919 3375 6957 3543
rect 6991 3375 7007 3543
rect 6919 3359 7007 3375
rect 6631 3285 6719 3301
rect 6631 3117 6647 3285
rect 6681 3117 6719 3285
rect 6631 3101 6719 3117
rect 6919 3285 7007 3301
rect 6919 3117 6957 3285
rect 6991 3117 7007 3285
rect 6919 3101 7007 3117
rect 7409 7871 7506 7887
rect 7409 7503 7425 7871
rect 7459 7503 7506 7871
rect 7409 7487 7506 7503
rect 7706 7871 7803 7887
rect 7706 7503 7753 7871
rect 7787 7503 7803 7871
rect 7706 7487 7803 7503
rect 7409 6581 7506 6597
rect 7409 6213 7425 6581
rect 7459 6213 7506 6581
rect 7409 6197 7506 6213
rect 7706 6581 7803 6597
rect 7706 6213 7753 6581
rect 7787 6213 7803 6581
rect 7706 6197 7803 6213
rect 17958 7207 18046 7223
rect 17958 6239 17974 7207
rect 18008 6239 18046 7207
rect 17958 6223 18046 6239
rect 18646 7207 18734 7223
rect 18646 6239 18684 7207
rect 18718 6239 18734 7207
rect 18646 6223 18734 6239
rect 19431 8866 21831 8882
rect 19431 8832 19447 8866
rect 21815 8832 21831 8866
rect 19431 8794 21831 8832
rect 21889 8866 24289 8882
rect 21889 8832 21905 8866
rect 24273 8832 24289 8866
rect 21889 8794 24289 8832
rect 19431 7556 21831 7594
rect 19431 7522 19447 7556
rect 21815 7522 21831 7556
rect 19431 7506 21831 7522
rect 21889 7556 24289 7594
rect 21889 7522 21905 7556
rect 24273 7522 24289 7556
rect 21889 7506 24289 7522
rect 19430 6991 21830 7007
rect 19430 6957 19446 6991
rect 21814 6957 21830 6991
rect 19430 6919 21830 6957
rect 21888 6991 24288 7007
rect 21888 6957 21904 6991
rect 24272 6957 24288 6991
rect 21888 6919 24288 6957
rect 19430 5681 21830 5719
rect 19430 5647 19446 5681
rect 21814 5647 21830 5681
rect 19430 5631 21830 5647
rect 21888 5681 24288 5719
rect 21888 5647 21904 5681
rect 24272 5647 24288 5681
rect 21888 5631 24288 5647
rect 7409 5291 7506 5307
rect 7409 4923 7425 5291
rect 7459 4923 7506 5291
rect 7409 4907 7506 4923
rect 7706 5291 7803 5307
rect 7706 4923 7753 5291
rect 7787 4923 7803 5291
rect 7706 4907 7803 4923
rect 7409 4001 7506 4017
rect 7409 3633 7425 4001
rect 7459 3633 7506 4001
rect 7409 3617 7506 3633
rect 7706 4001 7803 4017
rect 7706 3633 7753 4001
rect 7787 3633 7803 4001
rect 7706 3617 7803 3633
rect 7409 3420 7506 3436
rect 7409 3052 7425 3420
rect 7459 3052 7506 3420
rect 7409 3036 7506 3052
rect 7706 3420 7803 3436
rect 7706 3052 7753 3420
rect 7787 3052 7803 3420
rect 7706 3036 7803 3052
<< polycont >>
rect 3728 30499 7296 30533
rect 7386 30499 10954 30533
rect 3728 30011 7296 30045
rect 7386 30011 10954 30045
rect 3728 29523 7296 29557
rect 7386 29523 10954 29557
rect 3465 26025 3499 26993
rect 4175 26025 4209 26993
rect 4938 28618 7306 28652
rect 7396 28618 9764 28652
rect 4938 27308 7306 27342
rect 7396 27308 9764 27342
rect 4937 26743 7305 26777
rect 7395 26743 9763 26777
rect 4937 25433 7305 25467
rect 7395 25433 9763 25467
rect 12200 32575 12548 32609
rect 12638 32575 12986 32609
rect 13076 32575 13424 32609
rect 13514 32575 13862 32609
rect 12200 29447 12548 29481
rect 12638 29447 12986 29481
rect 13076 29447 13424 29481
rect 13514 29447 13862 29481
rect 12200 28598 12548 28632
rect 12638 28598 12986 28632
rect 13076 28598 13424 28632
rect 13514 28598 13862 28632
rect 12200 25470 12548 25504
rect 12638 25470 12986 25504
rect 13076 25470 13424 25504
rect 13514 25470 13862 25504
rect 17029 27044 17357 27078
rect 17447 27044 17775 27078
rect 17865 27044 18193 27078
rect 18283 27044 18611 27078
rect 17029 25516 17357 25550
rect 17447 25516 17775 25550
rect 17865 25516 18193 25550
rect 18283 25516 18611 25550
rect 21122 27589 22090 27623
rect 22180 27589 23148 27623
rect 23238 27589 24206 27623
rect 24296 27589 25264 27623
rect 21122 26961 22090 26995
rect 22180 26961 23148 26995
rect 23238 26961 24206 26995
rect 24296 26961 25264 26995
rect 21122 26427 22090 26461
rect 22180 26427 23148 26461
rect 23238 26427 24206 26461
rect 24296 26427 25264 26461
rect 21122 25799 22090 25833
rect 22180 25799 23148 25833
rect 23238 25799 24206 25833
rect 24296 25799 25264 25833
rect 12210 24563 14058 24597
rect 14148 24563 15996 24597
rect 16086 24563 17934 24597
rect 18024 24563 19872 24597
rect 12210 24153 14058 24187
rect 14148 24153 15996 24187
rect 16086 24153 17934 24187
rect 18024 24153 19872 24187
rect 12210 23743 14058 23777
rect 14148 23743 15996 23777
rect 16086 23743 17934 23777
rect 18024 23743 19872 23777
rect 22307 25133 22675 25167
rect 22765 25133 23133 25167
rect 23223 25133 23591 25167
rect 23681 25133 24049 25167
rect 22307 24423 22675 24457
rect 22765 24423 23133 24457
rect 23223 24423 23591 24457
rect 23681 24423 24049 24457
rect 22307 23926 22675 23960
rect 22765 23926 23133 23960
rect 23223 23926 23591 23960
rect 23681 23926 24049 23960
rect 22307 23216 22675 23250
rect 22765 23216 23133 23250
rect 23223 23216 23591 23250
rect 23681 23216 24049 23250
rect 25455 25024 25493 25058
rect 25455 24376 25493 24410
rect 25811 25024 25849 25058
rect 25811 24376 25849 24410
rect 25477 24010 25511 24044
rect 25833 24010 25867 24044
rect 25477 23700 25511 23734
rect 25833 23700 25867 23734
rect 12394 21340 12428 21508
rect 13304 21340 13338 21508
rect 13875 21340 13909 21508
rect 14785 21340 14819 21508
rect 12394 21082 12428 21250
rect 13304 21082 13338 21250
rect 13875 21082 13909 21250
rect 14785 21082 14819 21250
rect 12394 20824 12428 20992
rect 13304 20824 13338 20992
rect 13875 20824 13909 20992
rect 14785 20824 14819 20992
rect 12394 20566 12428 20734
rect 13304 20566 13338 20734
rect 13875 20566 13909 20734
rect 14785 20566 14819 20734
rect 12394 20308 12428 20476
rect 13304 20308 13338 20476
rect 13875 20308 13909 20476
rect 14785 20308 14819 20476
rect 12394 20050 12428 20218
rect 13304 20050 13338 20218
rect 13875 20050 13909 20218
rect 14785 20050 14819 20218
rect 12394 19792 12428 19960
rect 13304 19792 13338 19960
rect 13875 19792 13909 19960
rect 14785 19792 14819 19960
rect 12394 19534 12428 19702
rect 13304 19534 13338 19702
rect 13875 19534 13909 19702
rect 14785 19534 14819 19702
rect 12394 19276 12428 19444
rect 13304 19276 13338 19444
rect 13875 19276 13909 19444
rect 14785 19276 14819 19444
rect 12394 19018 12428 19186
rect 13304 19018 13338 19186
rect 13875 19018 13909 19186
rect 14785 19018 14819 19186
rect 12394 18760 12428 18928
rect 13304 18760 13338 18928
rect 13875 18760 13909 18928
rect 14785 18760 14819 18928
rect 12394 18502 12428 18670
rect 13304 18502 13338 18670
rect 13875 18502 13909 18670
rect 14785 18502 14819 18670
rect 12394 18244 12428 18412
rect 13304 18244 13338 18412
rect 13875 18244 13909 18412
rect 14785 18244 14819 18412
rect 12394 17986 12428 18154
rect 13304 17986 13338 18154
rect 13875 17986 13909 18154
rect 14785 17986 14819 18154
rect 12394 17728 12428 17896
rect 13304 17728 13338 17896
rect 13875 17728 13909 17896
rect 14785 17728 14819 17896
rect 12394 17470 12428 17638
rect 13304 17470 13338 17638
rect 13875 17470 13909 17638
rect 14785 17470 14819 17638
rect 12394 17212 12428 17380
rect 13304 17212 13338 17380
rect 13875 17212 13909 17380
rect 14785 17212 14819 17380
rect 12394 16954 12428 17122
rect 13304 16954 13338 17122
rect 13875 16954 13909 17122
rect 14785 16954 14819 17122
rect 12394 16696 12428 16864
rect 13304 16696 13338 16864
rect 13875 16696 13909 16864
rect 14785 16696 14819 16864
rect 12394 16438 12428 16606
rect 13304 16438 13338 16606
rect 13875 16438 13909 16606
rect 14785 16438 14819 16606
rect 12394 16180 12428 16348
rect 13304 16180 13338 16348
rect 13875 16180 13909 16348
rect 14785 16180 14819 16348
rect 12394 15922 12428 16090
rect 13304 15922 13338 16090
rect 13875 15922 13909 16090
rect 14785 15922 14819 16090
rect 12394 15664 12428 15832
rect 13304 15664 13338 15832
rect 13875 15664 13909 15832
rect 14785 15664 14819 15832
rect 12394 15406 12428 15574
rect 13304 15406 13338 15574
rect 13875 15406 13909 15574
rect 14785 15406 14819 15574
rect 16012 22145 16046 22313
rect 16322 22145 16356 22313
rect 16012 21887 16046 22055
rect 16322 21887 16356 22055
rect 16012 21629 16046 21797
rect 16322 21629 16356 21797
rect 16012 21371 16046 21539
rect 16322 21371 16356 21539
rect 16012 21113 16046 21281
rect 16322 21113 16356 21281
rect 16012 20855 16046 21023
rect 16322 20855 16356 21023
rect 16012 20597 16046 20765
rect 16322 20597 16356 20765
rect 16012 20339 16046 20507
rect 16322 20339 16356 20507
rect 16012 20081 16046 20249
rect 16322 20081 16356 20249
rect 16012 19823 16046 19991
rect 16322 19823 16356 19991
rect 16012 19565 16046 19733
rect 16322 19565 16356 19733
rect 16012 19307 16046 19475
rect 16322 19307 16356 19475
rect 16012 19049 16046 19217
rect 16322 19049 16356 19217
rect 16012 18791 16046 18959
rect 16322 18791 16356 18959
rect 16012 18533 16046 18701
rect 16322 18533 16356 18701
rect 16012 18275 16046 18443
rect 16322 18275 16356 18443
rect 16012 18017 16046 18185
rect 16322 18017 16356 18185
rect 16012 17759 16046 17927
rect 16322 17759 16356 17927
rect 16012 17501 16046 17669
rect 16322 17501 16356 17669
rect 16012 17243 16046 17411
rect 16322 17243 16356 17411
rect 16790 22010 16824 22378
rect 17118 22010 17152 22378
rect 16790 21429 16824 21797
rect 17118 21429 17152 21797
rect 22582 22420 22616 22688
rect 23792 22420 23826 22688
rect 22582 22062 22616 22330
rect 23792 22062 23826 22330
rect 16790 20139 16824 20507
rect 17118 20139 17152 20507
rect 16790 18849 16824 19217
rect 17118 18849 17152 19217
rect 16790 17559 16824 17927
rect 17118 17559 17152 17927
rect 16790 16671 16824 16839
rect 17118 16671 17152 16839
rect 16790 16413 16824 16581
rect 17118 16413 17152 16581
rect 16790 15746 16824 16114
rect 17018 15746 17052 16114
rect 16790 15288 16824 15656
rect 17018 15288 17052 15656
rect 3029 9955 3063 10123
rect 3939 9955 3973 10123
rect 4510 9955 4544 10123
rect 5420 9955 5454 10123
rect 3029 9697 3063 9865
rect 3939 9697 3973 9865
rect 4510 9697 4544 9865
rect 5420 9697 5454 9865
rect 3029 9439 3063 9607
rect 3939 9439 3973 9607
rect 4510 9439 4544 9607
rect 5420 9439 5454 9607
rect 3029 9181 3063 9349
rect 3939 9181 3973 9349
rect 4510 9181 4544 9349
rect 5420 9181 5454 9349
rect 3029 8923 3063 9091
rect 3939 8923 3973 9091
rect 4510 8923 4544 9091
rect 5420 8923 5454 9091
rect 3029 8665 3063 8833
rect 3939 8665 3973 8833
rect 4510 8665 4544 8833
rect 5420 8665 5454 8833
rect 3029 8407 3063 8575
rect 3939 8407 3973 8575
rect 4510 8407 4544 8575
rect 5420 8407 5454 8575
rect 3029 8149 3063 8317
rect 3939 8149 3973 8317
rect 4510 8149 4544 8317
rect 5420 8149 5454 8317
rect 3029 7891 3063 8059
rect 3939 7891 3973 8059
rect 4510 7891 4544 8059
rect 5420 7891 5454 8059
rect 3029 7633 3063 7801
rect 3939 7633 3973 7801
rect 4510 7633 4544 7801
rect 5420 7633 5454 7801
rect 3029 7375 3063 7543
rect 3939 7375 3973 7543
rect 4510 7375 4544 7543
rect 5420 7375 5454 7543
rect 3029 7117 3063 7285
rect 3939 7117 3973 7285
rect 4510 7117 4544 7285
rect 5420 7117 5454 7285
rect 3029 6859 3063 7027
rect 3939 6859 3973 7027
rect 4510 6859 4544 7027
rect 5420 6859 5454 7027
rect 3029 6601 3063 6769
rect 3939 6601 3973 6769
rect 4510 6601 4544 6769
rect 5420 6601 5454 6769
rect 3029 6343 3063 6511
rect 3939 6343 3973 6511
rect 4510 6343 4544 6511
rect 5420 6343 5454 6511
rect 3029 6085 3063 6253
rect 3939 6085 3973 6253
rect 4510 6085 4544 6253
rect 5420 6085 5454 6253
rect 3029 5827 3063 5995
rect 3939 5827 3973 5995
rect 4510 5827 4544 5995
rect 5420 5827 5454 5995
rect 3029 5569 3063 5737
rect 3939 5569 3973 5737
rect 4510 5569 4544 5737
rect 5420 5569 5454 5737
rect 3029 5311 3063 5479
rect 3939 5311 3973 5479
rect 4510 5311 4544 5479
rect 5420 5311 5454 5479
rect 3029 5053 3063 5221
rect 3939 5053 3973 5221
rect 4510 5053 4544 5221
rect 5420 5053 5454 5221
rect 3029 4795 3063 4963
rect 3939 4795 3973 4963
rect 4510 4795 4544 4963
rect 5420 4795 5454 4963
rect 3029 4537 3063 4705
rect 3939 4537 3973 4705
rect 4510 4537 4544 4705
rect 5420 4537 5454 4705
rect 3029 4279 3063 4447
rect 3939 4279 3973 4447
rect 4510 4279 4544 4447
rect 5420 4279 5454 4447
rect 3029 4021 3063 4189
rect 3939 4021 3973 4189
rect 4510 4021 4544 4189
rect 5420 4021 5454 4189
rect 7425 9873 7459 10241
rect 7653 9873 7687 10241
rect 7425 9415 7459 9783
rect 7653 9415 7687 9783
rect 7425 8948 7459 9116
rect 7753 8948 7787 9116
rect 7425 8690 7459 8858
rect 7753 8690 7787 8858
rect 18237 10713 21805 10747
rect 21895 10713 25463 10747
rect 18237 10225 21805 10259
rect 21895 10225 25463 10259
rect 18237 9737 21805 9771
rect 21895 9737 25463 9771
rect 6647 8019 6681 8187
rect 6957 8019 6991 8187
rect 6647 7761 6681 7929
rect 6957 7761 6991 7929
rect 6647 7503 6681 7671
rect 6957 7503 6991 7671
rect 6647 7245 6681 7413
rect 6957 7245 6991 7413
rect 6647 6987 6681 7155
rect 6957 6987 6991 7155
rect 6647 6729 6681 6897
rect 6957 6729 6991 6897
rect 6647 6471 6681 6639
rect 6957 6471 6991 6639
rect 6647 6213 6681 6381
rect 6957 6213 6991 6381
rect 6647 5955 6681 6123
rect 6957 5955 6991 6123
rect 6647 5697 6681 5865
rect 6957 5697 6991 5865
rect 6647 5439 6681 5607
rect 6957 5439 6991 5607
rect 6647 5181 6681 5349
rect 6957 5181 6991 5349
rect 6647 4923 6681 5091
rect 6957 4923 6991 5091
rect 6647 4665 6681 4833
rect 6957 4665 6991 4833
rect 6647 4407 6681 4575
rect 6957 4407 6991 4575
rect 6647 4149 6681 4317
rect 6957 4149 6991 4317
rect 6647 3891 6681 4059
rect 6957 3891 6991 4059
rect 6647 3633 6681 3801
rect 6957 3633 6991 3801
rect 6647 3375 6681 3543
rect 6957 3375 6991 3543
rect 6647 3117 6681 3285
rect 6957 3117 6991 3285
rect 7425 7503 7459 7871
rect 7753 7503 7787 7871
rect 7425 6213 7459 6581
rect 7753 6213 7787 6581
rect 17974 6239 18008 7207
rect 18684 6239 18718 7207
rect 19447 8832 21815 8866
rect 21905 8832 24273 8866
rect 19447 7522 21815 7556
rect 21905 7522 24273 7556
rect 19446 6957 21814 6991
rect 21904 6957 24272 6991
rect 19446 5647 21814 5681
rect 21904 5647 24272 5681
rect 7425 4923 7459 5291
rect 7753 4923 7787 5291
rect 7425 3633 7459 4001
rect 7753 3633 7787 4001
rect 7425 3052 7459 3420
rect 7753 3052 7787 3420
<< xpolycontact >>
rect 24889 22946 25321 23016
rect 25529 22946 25961 23016
<< xpolyres >>
rect 25321 22946 25529 23016
<< locali >>
rect 11766 33012 14431 33025
rect 3217 30890 11393 30926
rect 3217 30801 3401 30890
rect 11199 30801 11393 30890
rect 3217 30745 11393 30801
rect 3217 30711 3469 30745
rect 11157 30711 11393 30745
rect 3217 30685 11393 30711
rect 3217 29429 3409 30685
rect 3443 30588 11183 30685
rect 3443 29429 3471 30588
rect 3712 30499 3728 30533
rect 7296 30499 7312 30533
rect 7370 30499 7386 30533
rect 10954 30499 10970 30533
rect 3666 30440 3700 30456
rect 3666 30088 3700 30104
rect 7324 30440 7358 30456
rect 7324 30088 7358 30104
rect 10982 30440 11016 30456
rect 10982 30088 11016 30104
rect 3712 30011 3728 30045
rect 7296 30011 7312 30045
rect 7370 30011 7386 30045
rect 10954 30011 10970 30045
rect 3666 29952 3700 29968
rect 3666 29600 3700 29616
rect 7324 29952 7358 29968
rect 7324 29600 7358 29616
rect 10982 29952 11016 29968
rect 10982 29600 11016 29616
rect 3712 29523 3728 29557
rect 7296 29523 7312 29557
rect 7370 29523 7386 29557
rect 10954 29523 10970 29557
rect 3217 29419 3471 29429
rect 11217 30588 11393 30685
rect 11217 29429 11392 30588
rect 11183 29419 11392 29429
rect 3217 29403 11392 29419
rect 3217 29369 3469 29403
rect 11157 29369 11392 29403
rect 3217 29286 11392 29369
rect 11766 29401 11800 33012
rect 14392 32809 14431 33012
rect 11965 32791 14240 32809
rect 11965 29401 12000 32791
rect 12184 32575 12200 32609
rect 12548 32575 12564 32609
rect 12622 32575 12638 32609
rect 12986 32575 13002 32609
rect 13060 32575 13076 32609
rect 13424 32575 13440 32609
rect 13498 32575 13514 32609
rect 13862 32575 13878 32609
rect 12138 32516 12172 32532
rect 12138 29524 12172 29540
rect 12576 32516 12610 32532
rect 12576 29524 12610 29540
rect 13014 32516 13048 32532
rect 13014 29524 13048 29540
rect 13452 32516 13486 32532
rect 13452 29524 13486 29540
rect 13890 32516 13924 32532
rect 13890 29524 13924 29540
rect 14115 32230 14240 32791
rect 14274 32230 14431 32809
rect 14115 29750 14180 32230
rect 14322 29750 14431 32230
rect 12184 29447 12200 29481
rect 12548 29447 12564 29481
rect 12622 29447 12638 29481
rect 12986 29447 13002 29481
rect 13060 29447 13076 29481
rect 13424 29447 13440 29481
rect 13498 29447 13514 29481
rect 13862 29447 13878 29481
rect 3218 28784 10367 28851
rect 3218 28750 4700 28784
rect 10001 28750 10367 28784
rect 3218 28724 10367 28750
rect 3218 27170 4640 28724
rect 3217 27169 4640 27170
rect 3217 27135 3459 27169
rect 4215 27135 4640 27169
rect 3217 27133 4640 27135
rect 3217 27073 3428 27133
rect 3217 25945 3363 27073
rect 3397 25945 3428 27073
rect 4269 27073 4640 27133
rect 3533 27021 3549 27055
rect 4125 27021 4141 27055
rect 3465 26993 3499 27009
rect 3465 26009 3499 26025
rect 4175 26993 4209 27009
rect 4175 26009 4209 26025
rect 3217 25887 3428 25945
rect 3533 25963 3549 25997
rect 4125 25963 4141 25997
rect 3533 25887 4141 25963
rect 4269 25945 4277 27073
rect 4311 25945 4640 27073
rect 4269 25887 4640 25945
rect 3217 25883 4640 25887
rect 3217 25849 3459 25883
rect 4215 25849 4640 25883
rect 3217 25657 4640 25849
rect 3215 25453 4640 25657
rect 3215 25359 3323 25453
rect 3876 25382 4640 25453
rect 4674 28711 10027 28724
rect 4674 25382 4694 28711
rect 4922 28618 4938 28652
rect 7306 28618 7322 28652
rect 7380 28618 7396 28652
rect 9764 28618 9780 28652
rect 4876 28568 4910 28584
rect 4876 27376 4910 27392
rect 7334 28568 7368 28584
rect 7334 27376 7368 27392
rect 9792 28568 9826 28584
rect 9792 27376 9826 27392
rect 4922 27308 4938 27342
rect 7306 27308 7322 27342
rect 7380 27308 7396 27342
rect 9764 27308 9780 27342
rect 4921 26743 4937 26777
rect 7305 26743 7321 26777
rect 7379 26743 7395 26777
rect 9763 26743 9779 26777
rect 4875 26693 4909 26709
rect 4875 25501 4909 25517
rect 7333 26693 7367 26709
rect 7333 25501 7367 25517
rect 9791 26693 9825 26709
rect 9791 25501 9825 25517
rect 4921 25433 4937 25467
rect 7305 25433 7321 25467
rect 7379 25433 7395 25467
rect 9763 25433 9779 25467
rect 3876 25377 4694 25382
rect 10017 25382 10027 28711
rect 10061 25382 10367 28724
rect 10017 25377 10367 25382
rect 3876 25359 10367 25377
rect 3215 25356 10367 25359
rect 3215 25322 4700 25356
rect 10001 25322 10367 25356
rect 3215 25218 10367 25322
rect 11766 28583 11874 29401
rect 11908 28583 12000 29401
rect 12184 28598 12200 28632
rect 12548 28598 12564 28632
rect 12622 28598 12638 28632
rect 12986 28598 13002 28632
rect 13060 28598 13076 28632
rect 13424 28598 13440 28632
rect 13498 28598 13514 28632
rect 13862 28598 13878 28632
rect 11766 25407 11817 28583
rect 11766 25231 11816 25407
rect 11965 25388 12000 28583
rect 12138 28539 12172 28555
rect 12138 25547 12172 25563
rect 12576 28539 12610 28555
rect 12576 25547 12610 25563
rect 13014 28539 13048 28555
rect 13014 25547 13048 25563
rect 13452 28539 13486 28555
rect 13452 25547 13486 25563
rect 13890 28539 13924 28555
rect 13890 25547 13924 25563
rect 14115 27997 14240 29750
rect 14274 27997 14431 29750
rect 14115 25517 14196 27997
rect 14338 27586 14431 27997
rect 20550 28158 25680 28530
rect 20550 28157 25403 28158
rect 20550 27792 20700 28157
rect 25662 27826 25680 28158
rect 20550 27680 20762 27792
rect 14338 27499 19171 27586
rect 19128 27498 19171 27499
rect 14338 27120 16600 27207
rect 14338 25517 14431 27120
rect 12184 25470 12200 25504
rect 12548 25470 12564 25504
rect 12622 25470 12638 25504
rect 12986 25470 13002 25504
rect 13060 25470 13076 25504
rect 13424 25470 13440 25504
rect 13498 25470 13514 25504
rect 13862 25470 13878 25504
rect 14115 25388 14240 25517
rect 11965 25374 14240 25388
rect 14274 25374 14431 25517
rect 14381 25250 14431 25374
rect 11766 25230 11929 25231
rect 14381 25230 14417 25250
rect 11766 25223 14417 25230
rect 3215 25129 3325 25218
rect 10259 25129 10367 25218
rect 16555 25217 16600 27120
rect 16833 27180 18851 27207
rect 16833 27146 16949 27180
rect 18691 27146 18851 27180
rect 16833 27120 18851 27146
rect 16833 27084 16897 27120
rect 16833 25510 16853 27084
rect 16887 25510 16897 27084
rect 18737 27084 18851 27120
rect 17013 27044 17029 27078
rect 17357 27044 17373 27078
rect 17431 27044 17447 27078
rect 17775 27044 17791 27078
rect 17849 27044 17865 27078
rect 18193 27044 18209 27078
rect 18267 27044 18283 27078
rect 18611 27044 18627 27078
rect 16967 26985 17001 27001
rect 16967 25593 17001 25609
rect 17385 26985 17419 27001
rect 17385 25593 17419 25609
rect 17803 26985 17837 27001
rect 17803 25593 17837 25609
rect 18221 26985 18255 27001
rect 18221 25593 18255 25609
rect 18639 26985 18673 27001
rect 18639 25593 18673 25609
rect 17013 25516 17029 25550
rect 17357 25516 17373 25550
rect 17431 25516 17447 25550
rect 17775 25516 17791 25550
rect 17849 25516 17865 25550
rect 18193 25516 18209 25550
rect 18267 25516 18283 25550
rect 18611 25516 18627 25550
rect 16833 25477 16897 25510
rect 18737 25510 18753 27084
rect 18787 25691 18851 27084
rect 19138 25691 19171 27498
rect 18787 25510 19171 25691
rect 18737 25477 19171 25510
rect 16833 25457 19171 25477
rect 20741 25500 20762 27680
rect 25504 27792 25546 27793
rect 20879 27680 25546 27792
rect 20879 25624 20921 27680
rect 21106 27589 21122 27623
rect 22090 27589 22106 27623
rect 22164 27589 22180 27623
rect 23148 27589 23164 27623
rect 23222 27589 23238 27623
rect 24206 27589 24222 27623
rect 24280 27589 24296 27623
rect 25264 27589 25280 27623
rect 21060 27530 21094 27546
rect 21060 27038 21094 27054
rect 22118 27530 22152 27546
rect 22118 27038 22152 27054
rect 23176 27530 23210 27546
rect 23176 27038 23210 27054
rect 24234 27530 24268 27546
rect 24234 27038 24268 27054
rect 25292 27530 25326 27546
rect 25292 27038 25326 27054
rect 21106 26961 21122 26995
rect 22090 26961 22106 26995
rect 22164 26961 22180 26995
rect 23148 26961 23164 26995
rect 23222 26961 23238 26995
rect 24206 26961 24222 26995
rect 24280 26961 24296 26995
rect 25264 26961 25280 26995
rect 25525 26979 25546 27680
rect 25662 27793 25683 27826
rect 25643 26979 25683 27793
rect 21106 26427 21122 26461
rect 22090 26427 22106 26461
rect 22164 26427 22180 26461
rect 23148 26427 23164 26461
rect 23222 26427 23238 26461
rect 24206 26427 24222 26461
rect 24280 26427 24296 26461
rect 25264 26427 25280 26461
rect 21060 26368 21094 26384
rect 21060 25876 21094 25892
rect 22118 26368 22152 26384
rect 22118 25876 22152 25892
rect 23176 26368 23210 26384
rect 23176 25876 23210 25892
rect 24234 26368 24268 26384
rect 24234 25876 24268 25892
rect 25292 26368 25326 26384
rect 25292 25876 25326 25892
rect 21106 25799 21122 25833
rect 22090 25799 22106 25833
rect 22164 25799 22180 25833
rect 23148 25799 23164 25833
rect 23222 25799 23238 25833
rect 24206 25799 24222 25833
rect 24280 25799 24296 25833
rect 25264 25799 25280 25833
rect 25525 25624 25567 26979
rect 20879 25590 25567 25624
rect 25311 25585 25567 25590
rect 25601 25585 25683 26979
rect 25311 25559 25683 25585
rect 25541 25548 25683 25559
rect 25541 25525 26070 25548
rect 20741 25493 20797 25500
rect 20741 25472 25207 25493
rect 20755 25466 25207 25472
rect 16833 25451 19175 25457
rect 16555 25215 16685 25217
rect 18748 25215 19175 25451
rect 22093 25360 24294 25385
rect 22093 25235 22120 25360
rect 24269 25263 24294 25360
rect 16555 25201 19175 25215
rect 3215 25067 10367 25129
rect 11862 24892 19698 24929
rect 11862 23392 11872 24892
rect 12019 24889 19698 24892
rect 19814 24889 20269 24929
rect 20155 24855 20269 24889
rect 19814 24829 20269 24855
rect 12019 24768 19698 24780
rect 19814 24768 20181 24829
rect 12019 24742 20181 24768
rect 12019 23664 12040 24742
rect 12194 24563 12210 24597
rect 14058 24563 14074 24597
rect 14132 24563 14148 24597
rect 15996 24563 16012 24597
rect 16070 24563 16086 24597
rect 17934 24563 17950 24597
rect 18008 24563 18024 24597
rect 19872 24563 19888 24597
rect 12148 24513 12182 24529
rect 12148 24221 12182 24237
rect 14086 24513 14120 24529
rect 14086 24221 14120 24237
rect 16024 24513 16058 24529
rect 16024 24221 16058 24237
rect 17962 24513 17996 24529
rect 17962 24221 17996 24237
rect 19900 24513 19934 24529
rect 19900 24221 19934 24237
rect 12194 24153 12210 24187
rect 14058 24153 14074 24187
rect 14132 24153 14148 24187
rect 15996 24153 16012 24187
rect 16070 24153 16086 24187
rect 17934 24153 17950 24187
rect 18008 24153 18024 24187
rect 19872 24153 19888 24187
rect 12148 24103 12182 24119
rect 12148 23811 12182 23827
rect 14086 24103 14120 24119
rect 14086 23811 14120 23827
rect 16024 24103 16058 24119
rect 16024 23811 16058 23827
rect 17962 24103 17996 24119
rect 17962 23811 17996 23827
rect 19900 24103 19934 24119
rect 19900 23811 19934 23827
rect 12194 23743 12210 23777
rect 14058 23743 14074 23777
rect 14132 23743 14148 23777
rect 15996 23743 16012 23777
rect 16070 23743 16086 23777
rect 17934 23743 17950 23777
rect 18008 23743 18024 23777
rect 19872 23743 19888 23777
rect 20100 23664 20181 24742
rect 12019 23606 20181 23664
rect 20215 23606 20269 24829
rect 12019 23590 20269 23606
rect 12113 23589 20269 23590
rect 19791 23580 20269 23589
rect 20155 23546 20269 23580
rect 19791 23392 20269 23546
rect 11862 23375 20269 23392
rect 11871 23374 20269 23375
rect 22100 24719 22120 25235
rect 22178 25235 24193 25257
rect 22178 24719 22193 25235
rect 22291 25133 22307 25167
rect 22675 25133 22691 25167
rect 22749 25133 22765 25167
rect 23133 25133 23149 25167
rect 23207 25133 23223 25167
rect 23591 25133 23607 25167
rect 23665 25133 23681 25167
rect 24049 25133 24065 25167
rect 22100 23683 22135 24719
rect 22169 23683 22193 24719
rect 22245 25083 22279 25099
rect 22245 24491 22279 24507
rect 22703 25083 22737 25099
rect 22703 24491 22737 24507
rect 23161 25083 23195 25099
rect 23161 24491 23195 24507
rect 23619 25083 23653 25099
rect 23619 24491 23653 24507
rect 24077 25083 24111 25099
rect 24077 24491 24111 24507
rect 22291 24423 22307 24457
rect 22675 24423 22691 24457
rect 22749 24423 22765 24457
rect 23133 24423 23149 24457
rect 23207 24423 23223 24457
rect 23591 24423 23607 24457
rect 23665 24423 23681 24457
rect 24049 24423 24065 24457
rect 22291 23926 22307 23960
rect 22675 23926 22691 23960
rect 22749 23926 22765 23960
rect 23133 23926 23149 23960
rect 23207 23926 23223 23960
rect 23591 23926 23607 23960
rect 23665 23926 23681 23960
rect 24049 23926 24065 23960
rect 22100 23153 22111 23683
rect 22054 23052 22111 23153
rect 22185 23153 22193 23683
rect 22245 23876 22279 23892
rect 22245 23284 22279 23300
rect 22703 23876 22737 23892
rect 22703 23284 22737 23300
rect 23161 23876 23195 23892
rect 23161 23284 23195 23300
rect 23619 23876 23653 23892
rect 23619 23284 23653 23300
rect 24077 23876 24111 23892
rect 24077 23284 24111 23300
rect 22291 23216 22307 23250
rect 22675 23216 22691 23250
rect 22749 23216 22765 23250
rect 23133 23216 23149 23250
rect 23207 23216 23223 23250
rect 23591 23216 23607 23250
rect 23665 23216 23681 23250
rect 24049 23216 24065 23250
rect 24180 23153 24193 25235
rect 22185 23107 24193 23153
rect 24269 23154 24302 25263
rect 25186 24334 25207 25466
rect 25311 25160 26070 25525
rect 25311 25126 25375 25160
rect 25573 25126 25731 25160
rect 25929 25126 26070 25160
rect 25311 25107 26070 25126
rect 25311 25064 25324 25107
rect 25313 24370 25324 25064
rect 25635 25064 25669 25107
rect 25439 25024 25455 25058
rect 25493 25024 25509 25058
rect 25393 24965 25427 24981
rect 25393 24453 25427 24469
rect 25521 24965 25555 24981
rect 25521 24453 25555 24469
rect 25439 24376 25455 24410
rect 25493 24376 25509 24410
rect 25311 24334 25324 24370
rect 25186 24308 25324 24334
rect 25987 25064 26070 25107
rect 25795 25024 25811 25058
rect 25849 25024 25865 25058
rect 25749 24965 25783 24981
rect 25749 24453 25783 24469
rect 25877 24965 25911 24981
rect 25877 24453 25911 24469
rect 25795 24376 25811 24410
rect 25849 24376 25865 24410
rect 25635 24308 25669 24370
rect 25987 24370 25991 25064
rect 26025 24370 26070 25064
rect 25987 24308 26070 24370
rect 25186 24274 25375 24308
rect 25573 24274 25731 24308
rect 25929 24274 26070 24308
rect 25186 24251 25324 24274
rect 25987 24265 26070 24274
rect 24588 24146 26122 24166
rect 24588 24112 25371 24146
rect 25970 24112 26122 24146
rect 24588 24088 26122 24112
rect 24588 24086 25363 24088
rect 24588 23646 25311 24086
rect 25345 23646 25363 24086
rect 25976 24086 26122 24088
rect 25461 24010 25477 24044
rect 25511 24010 25527 24044
rect 25817 24010 25833 24044
rect 25867 24010 25883 24044
rect 25433 23960 25467 23976
rect 25433 23768 25467 23784
rect 25521 23960 25555 23976
rect 25521 23768 25555 23784
rect 25789 23960 25823 23976
rect 25789 23768 25823 23784
rect 25877 23960 25911 23976
rect 25877 23768 25911 23784
rect 25461 23700 25477 23734
rect 25511 23700 25527 23734
rect 25817 23700 25833 23734
rect 25867 23700 25883 23734
rect 24588 23637 25363 23646
rect 25976 23646 25996 24086
rect 26030 23646 26122 24086
rect 25976 23637 26122 23646
rect 24588 23620 26122 23637
rect 24588 23586 25371 23620
rect 25970 23586 26122 23620
rect 24588 23500 26122 23586
rect 24588 23154 24611 23500
rect 25989 23228 26122 23500
rect 22185 23073 22195 23107
rect 24177 23073 24193 23107
rect 22185 23052 24193 23073
rect 24269 23052 24611 23154
rect 24731 23146 26122 23228
rect 24731 23112 24855 23146
rect 25995 23112 26122 23146
rect 24731 23090 26122 23112
rect 22054 22815 22066 23052
rect 24731 23050 24793 23090
rect 24731 22912 24759 23050
rect 26051 23050 26122 23090
rect 24731 22882 24793 22912
rect 16672 22598 17216 22599
rect 15708 22542 16598 22589
rect 15708 22508 15898 22542
rect 16480 22508 16598 22542
rect 15708 22482 16598 22508
rect 15708 22467 15838 22482
rect 15872 22467 16506 22482
rect 15708 21740 15736 22467
rect 15155 21737 15736 21740
rect 11975 21714 15736 21737
rect 11975 21700 12250 21714
rect 11975 15122 12053 21700
rect 12227 21680 12250 21700
rect 14959 21680 15736 21714
rect 12227 21656 15736 21680
rect 12227 21654 14994 21656
rect 12227 21621 14985 21654
rect 12227 15198 12336 21621
rect 12462 21536 12478 21570
rect 13254 21536 13270 21570
rect 13943 21536 13959 21570
rect 14735 21536 14751 21570
rect 12394 21508 12428 21524
rect 12394 21324 12428 21340
rect 13304 21508 13338 21524
rect 13304 21324 13338 21340
rect 13875 21508 13909 21524
rect 13875 21324 13909 21340
rect 14785 21508 14819 21524
rect 14785 21324 14819 21340
rect 12462 21278 12478 21312
rect 13254 21278 13270 21312
rect 13943 21278 13959 21312
rect 14735 21278 14751 21312
rect 12394 21250 12428 21266
rect 12394 21066 12428 21082
rect 13304 21250 13338 21266
rect 13304 21066 13338 21082
rect 13875 21250 13909 21266
rect 13875 21066 13909 21082
rect 14785 21250 14819 21266
rect 14785 21066 14819 21082
rect 12462 21020 12478 21054
rect 13254 21020 13270 21054
rect 13943 21020 13959 21054
rect 14735 21020 14751 21054
rect 12394 20992 12428 21008
rect 12394 20808 12428 20824
rect 13304 20992 13338 21008
rect 13304 20808 13338 20824
rect 13875 20992 13909 21008
rect 13875 20808 13909 20824
rect 14785 20992 14819 21008
rect 14785 20808 14819 20824
rect 12462 20762 12478 20796
rect 13254 20762 13270 20796
rect 13943 20762 13959 20796
rect 14735 20762 14751 20796
rect 12394 20734 12428 20750
rect 12394 20550 12428 20566
rect 13304 20734 13338 20750
rect 13304 20550 13338 20566
rect 13875 20734 13909 20750
rect 13875 20550 13909 20566
rect 14785 20734 14819 20750
rect 14785 20550 14819 20566
rect 12462 20504 12478 20538
rect 13254 20504 13270 20538
rect 13943 20504 13959 20538
rect 14735 20504 14751 20538
rect 12394 20476 12428 20492
rect 12394 20292 12428 20308
rect 13304 20476 13338 20492
rect 13304 20292 13338 20308
rect 13875 20476 13909 20492
rect 13875 20292 13909 20308
rect 14785 20476 14819 20492
rect 14785 20292 14819 20308
rect 12462 20246 12478 20280
rect 13254 20246 13270 20280
rect 13943 20246 13959 20280
rect 14735 20246 14751 20280
rect 12394 20218 12428 20234
rect 12394 20034 12428 20050
rect 13304 20218 13338 20234
rect 13304 20034 13338 20050
rect 13875 20218 13909 20234
rect 13875 20034 13909 20050
rect 14785 20218 14819 20234
rect 14785 20034 14819 20050
rect 12462 19988 12478 20022
rect 13254 19988 13270 20022
rect 13943 19988 13959 20022
rect 14735 19988 14751 20022
rect 12394 19960 12428 19976
rect 12394 19776 12428 19792
rect 13304 19960 13338 19976
rect 13304 19776 13338 19792
rect 13875 19960 13909 19976
rect 13875 19776 13909 19792
rect 14785 19960 14819 19976
rect 14785 19776 14819 19792
rect 12462 19730 12478 19764
rect 13254 19730 13270 19764
rect 13943 19730 13959 19764
rect 14735 19730 14751 19764
rect 12394 19702 12428 19718
rect 12394 19518 12428 19534
rect 13304 19702 13338 19718
rect 13304 19518 13338 19534
rect 13875 19702 13909 19718
rect 13875 19518 13909 19534
rect 14785 19702 14819 19718
rect 14785 19518 14819 19534
rect 12462 19472 12478 19506
rect 13254 19472 13270 19506
rect 13943 19472 13959 19506
rect 14735 19472 14751 19506
rect 12394 19444 12428 19460
rect 12394 19260 12428 19276
rect 13304 19444 13338 19460
rect 13304 19260 13338 19276
rect 13875 19444 13909 19460
rect 13875 19260 13909 19276
rect 14785 19444 14819 19460
rect 14785 19260 14819 19276
rect 12462 19214 12478 19248
rect 13254 19214 13270 19248
rect 13943 19214 13959 19248
rect 14735 19214 14751 19248
rect 12394 19186 12428 19202
rect 12394 19002 12428 19018
rect 13304 19186 13338 19202
rect 13304 19002 13338 19018
rect 13875 19186 13909 19202
rect 13875 19002 13909 19018
rect 14785 19186 14819 19202
rect 14785 19002 14819 19018
rect 12462 18956 12478 18990
rect 13254 18956 13270 18990
rect 13943 18956 13959 18990
rect 14735 18956 14751 18990
rect 12394 18928 12428 18944
rect 12394 18744 12428 18760
rect 13304 18928 13338 18944
rect 13304 18744 13338 18760
rect 13875 18928 13909 18944
rect 13875 18744 13909 18760
rect 14785 18928 14819 18944
rect 14785 18744 14819 18760
rect 12462 18698 12478 18732
rect 13254 18698 13270 18732
rect 13943 18698 13959 18732
rect 14735 18698 14751 18732
rect 12394 18670 12428 18686
rect 12394 18486 12428 18502
rect 13304 18670 13338 18686
rect 13304 18486 13338 18502
rect 13875 18670 13909 18686
rect 13875 18486 13909 18502
rect 14785 18670 14819 18686
rect 14785 18486 14819 18502
rect 12462 18440 12478 18474
rect 13254 18440 13270 18474
rect 13943 18440 13959 18474
rect 14735 18440 14751 18474
rect 12394 18412 12428 18428
rect 12394 18228 12428 18244
rect 13304 18412 13338 18428
rect 13304 18228 13338 18244
rect 13875 18412 13909 18428
rect 13875 18228 13909 18244
rect 14785 18412 14819 18428
rect 14785 18228 14819 18244
rect 12462 18182 12478 18216
rect 13254 18182 13270 18216
rect 13943 18182 13959 18216
rect 14735 18182 14751 18216
rect 12394 18154 12428 18170
rect 12394 17970 12428 17986
rect 13304 18154 13338 18170
rect 13304 17970 13338 17986
rect 13875 18154 13909 18170
rect 13875 17970 13909 17986
rect 14785 18154 14819 18170
rect 14785 17970 14819 17986
rect 12462 17924 12478 17958
rect 13254 17924 13270 17958
rect 13943 17924 13959 17958
rect 14735 17924 14751 17958
rect 12394 17896 12428 17912
rect 12394 17712 12428 17728
rect 13304 17896 13338 17912
rect 13304 17712 13338 17728
rect 13875 17896 13909 17912
rect 13875 17712 13909 17728
rect 14785 17896 14819 17912
rect 14785 17712 14819 17728
rect 12462 17666 12478 17700
rect 13254 17666 13270 17700
rect 13943 17666 13959 17700
rect 14735 17666 14751 17700
rect 12394 17638 12428 17654
rect 12394 17454 12428 17470
rect 13304 17638 13338 17654
rect 13304 17454 13338 17470
rect 13875 17638 13909 17654
rect 13875 17454 13909 17470
rect 14785 17638 14819 17654
rect 14785 17454 14819 17470
rect 12462 17408 12478 17442
rect 13254 17408 13270 17442
rect 13943 17408 13959 17442
rect 14735 17408 14751 17442
rect 12394 17380 12428 17396
rect 12394 17196 12428 17212
rect 13304 17380 13338 17396
rect 13304 17196 13338 17212
rect 13875 17380 13909 17396
rect 13875 17196 13909 17212
rect 14785 17380 14819 17396
rect 14785 17196 14819 17212
rect 12462 17150 12478 17184
rect 13254 17150 13270 17184
rect 13943 17150 13959 17184
rect 14735 17150 14751 17184
rect 12394 17122 12428 17138
rect 12394 16938 12428 16954
rect 13304 17122 13338 17138
rect 13304 16938 13338 16954
rect 13875 17122 13909 17138
rect 13875 16938 13909 16954
rect 14785 17122 14819 17138
rect 14785 16938 14819 16954
rect 12462 16892 12478 16926
rect 13254 16892 13270 16926
rect 13943 16892 13959 16926
rect 14735 16892 14751 16926
rect 12394 16864 12428 16880
rect 12394 16680 12428 16696
rect 13304 16864 13338 16880
rect 13304 16680 13338 16696
rect 13875 16864 13909 16880
rect 13875 16680 13909 16696
rect 14785 16864 14819 16880
rect 14785 16680 14819 16696
rect 12462 16634 12478 16668
rect 13254 16634 13270 16668
rect 13943 16634 13959 16668
rect 14735 16634 14751 16668
rect 12394 16606 12428 16622
rect 12394 16422 12428 16438
rect 13304 16606 13338 16622
rect 13304 16422 13338 16438
rect 13875 16606 13909 16622
rect 13875 16422 13909 16438
rect 14785 16606 14819 16622
rect 14785 16422 14819 16438
rect 12462 16376 12478 16410
rect 13254 16376 13270 16410
rect 13943 16376 13959 16410
rect 14735 16376 14751 16410
rect 12394 16348 12428 16364
rect 12394 16164 12428 16180
rect 13304 16348 13338 16364
rect 13304 16164 13338 16180
rect 13875 16348 13909 16364
rect 13875 16164 13909 16180
rect 14785 16348 14819 16364
rect 14785 16164 14819 16180
rect 12462 16118 12478 16152
rect 13254 16118 13270 16152
rect 13943 16118 13959 16152
rect 14735 16118 14751 16152
rect 12394 16090 12428 16106
rect 12394 15906 12428 15922
rect 13304 16090 13338 16106
rect 13304 15906 13338 15922
rect 13875 16090 13909 16106
rect 13875 15906 13909 15922
rect 14785 16090 14819 16106
rect 14785 15906 14819 15922
rect 12462 15860 12478 15894
rect 13254 15860 13270 15894
rect 13943 15860 13959 15894
rect 14735 15860 14751 15894
rect 12394 15832 12428 15848
rect 12394 15648 12428 15664
rect 13304 15832 13338 15848
rect 13304 15648 13338 15664
rect 13875 15832 13909 15848
rect 13875 15648 13909 15664
rect 14785 15832 14819 15848
rect 14785 15648 14819 15664
rect 12462 15602 12478 15636
rect 13254 15602 13270 15636
rect 13943 15602 13959 15636
rect 14735 15602 14751 15636
rect 12394 15574 12428 15590
rect 12394 15390 12428 15406
rect 13304 15574 13338 15590
rect 13304 15390 13338 15406
rect 13875 15574 13909 15590
rect 13875 15390 13909 15406
rect 14785 15574 14819 15590
rect 14785 15390 14819 15406
rect 12462 15344 12478 15378
rect 13254 15344 13270 15378
rect 13943 15344 13959 15378
rect 14735 15344 14751 15378
rect 14942 15358 14985 21621
rect 14949 15198 14985 15358
rect 15106 17060 15736 21656
rect 15927 22466 16506 22467
rect 15927 17090 15964 22466
rect 16080 22341 16096 22375
rect 16272 22341 16288 22375
rect 16012 22313 16046 22329
rect 16012 22129 16046 22145
rect 16322 22313 16356 22329
rect 16322 22129 16356 22145
rect 16080 22083 16096 22117
rect 16272 22083 16288 22117
rect 16012 22055 16046 22071
rect 16012 21871 16046 21887
rect 16322 22055 16356 22071
rect 16322 21871 16356 21887
rect 16080 21825 16096 21859
rect 16272 21825 16288 21859
rect 16012 21797 16046 21813
rect 16012 21613 16046 21629
rect 16322 21797 16356 21813
rect 16322 21613 16356 21629
rect 16080 21567 16096 21601
rect 16272 21567 16288 21601
rect 16012 21539 16046 21555
rect 16012 21355 16046 21371
rect 16322 21539 16356 21555
rect 16322 21355 16356 21371
rect 16080 21309 16096 21343
rect 16272 21309 16288 21343
rect 16012 21281 16046 21297
rect 16012 21097 16046 21113
rect 16322 21281 16356 21297
rect 16322 21097 16356 21113
rect 16080 21051 16096 21085
rect 16272 21051 16288 21085
rect 16012 21023 16046 21039
rect 16012 20839 16046 20855
rect 16322 21023 16356 21039
rect 16322 20839 16356 20855
rect 16080 20793 16096 20827
rect 16272 20793 16288 20827
rect 16012 20765 16046 20781
rect 16012 20581 16046 20597
rect 16322 20765 16356 20781
rect 16322 20581 16356 20597
rect 16080 20535 16096 20569
rect 16272 20535 16288 20569
rect 16012 20507 16046 20523
rect 16012 20323 16046 20339
rect 16322 20507 16356 20523
rect 16322 20323 16356 20339
rect 16080 20277 16096 20311
rect 16272 20277 16288 20311
rect 16012 20249 16046 20265
rect 16012 20065 16046 20081
rect 16322 20249 16356 20265
rect 16322 20065 16356 20081
rect 16080 20019 16096 20053
rect 16272 20019 16288 20053
rect 16012 19991 16046 20007
rect 16012 19807 16046 19823
rect 16322 19991 16356 20007
rect 16322 19807 16356 19823
rect 16080 19761 16096 19795
rect 16272 19761 16288 19795
rect 16012 19733 16046 19749
rect 16012 19549 16046 19565
rect 16322 19733 16356 19749
rect 16322 19549 16356 19565
rect 16080 19503 16096 19537
rect 16272 19503 16288 19537
rect 16012 19475 16046 19491
rect 16012 19291 16046 19307
rect 16322 19475 16356 19491
rect 16322 19291 16356 19307
rect 16080 19245 16096 19279
rect 16272 19245 16288 19279
rect 16012 19217 16046 19233
rect 16012 19033 16046 19049
rect 16322 19217 16356 19233
rect 16322 19033 16356 19049
rect 16080 18987 16096 19021
rect 16272 18987 16288 19021
rect 16012 18959 16046 18975
rect 16012 18775 16046 18791
rect 16322 18959 16356 18975
rect 16322 18775 16356 18791
rect 16080 18729 16096 18763
rect 16272 18729 16288 18763
rect 16012 18701 16046 18717
rect 16012 18517 16046 18533
rect 16322 18701 16356 18717
rect 16322 18517 16356 18533
rect 16080 18471 16096 18505
rect 16272 18471 16288 18505
rect 16012 18443 16046 18459
rect 16012 18259 16046 18275
rect 16322 18443 16356 18459
rect 16322 18259 16356 18275
rect 16080 18213 16096 18247
rect 16272 18213 16288 18247
rect 16012 18185 16046 18201
rect 16012 18001 16046 18017
rect 16322 18185 16356 18201
rect 16322 18001 16356 18017
rect 16080 17955 16096 17989
rect 16272 17955 16288 17989
rect 16012 17927 16046 17943
rect 16012 17743 16046 17759
rect 16322 17927 16356 17943
rect 16322 17743 16356 17759
rect 16080 17697 16096 17731
rect 16272 17697 16288 17731
rect 16012 17669 16046 17685
rect 16012 17485 16046 17501
rect 16322 17669 16356 17685
rect 16322 17485 16356 17501
rect 16080 17439 16096 17473
rect 16272 17439 16288 17473
rect 16012 17411 16046 17427
rect 16012 17227 16046 17243
rect 16322 17411 16356 17427
rect 16322 17227 16356 17243
rect 16080 17181 16096 17215
rect 16272 17181 16288 17215
rect 16459 17090 16506 22466
rect 15927 17074 16506 17090
rect 16540 17074 16598 22482
rect 16672 22550 17624 22598
rect 16672 22516 16772 22550
rect 17196 22516 17624 22550
rect 16672 22495 17624 22516
rect 16672 22490 16751 22495
rect 16672 21326 16712 22490
rect 16746 21326 16751 22490
rect 17200 22490 17624 22495
rect 16867 22406 16883 22440
rect 17059 22406 17075 22440
rect 16790 22378 16824 22394
rect 16790 21994 16824 22010
rect 17118 22378 17152 22394
rect 17118 21994 17152 22010
rect 16867 21948 16883 21982
rect 17059 21948 17075 21982
rect 16867 21825 16883 21859
rect 17059 21825 17075 21859
rect 16790 21797 16824 21813
rect 16790 21413 16824 21429
rect 17118 21797 17152 21813
rect 17118 21413 17152 21429
rect 16867 21367 16883 21401
rect 17059 21367 17075 21401
rect 16672 21312 16751 21326
rect 17200 21326 17222 22490
rect 17256 22485 17624 22490
rect 17256 21326 17330 22485
rect 17200 21312 17330 21326
rect 16672 21300 17330 21312
rect 16672 21266 16772 21300
rect 17196 21266 17330 21300
rect 16672 21229 17330 21266
rect 16674 21227 17330 21229
rect 16838 20719 17330 21227
rect 16663 20683 17330 20719
rect 16663 20649 16784 20683
rect 17158 20649 17330 20683
rect 16663 20623 17330 20649
rect 16663 20587 16746 20623
rect 17199 20622 17330 20623
rect 16663 20059 16688 20587
rect 16722 20059 16746 20587
rect 17200 20587 17330 20622
rect 16867 20535 16883 20569
rect 17059 20535 17075 20569
rect 16790 20507 16824 20523
rect 16790 20123 16824 20139
rect 17118 20507 17152 20523
rect 17118 20123 17152 20139
rect 17200 20122 17220 20587
rect 16867 20077 16883 20111
rect 17059 20077 17075 20111
rect 16663 20026 16746 20059
rect 17199 20059 17220 20122
rect 17254 20059 17330 20587
rect 17199 20026 17330 20059
rect 16663 19997 17330 20026
rect 16663 19963 16784 19997
rect 17158 19963 17330 19997
rect 16663 19935 17330 19963
rect 16838 19429 17330 19935
rect 16672 19393 17330 19429
rect 16672 19359 16784 19393
rect 17158 19359 17330 19393
rect 16672 19349 17330 19359
rect 16672 19297 16748 19349
rect 16672 18769 16688 19297
rect 16722 18769 16748 19297
rect 17200 19297 17330 19349
rect 16867 19245 16883 19279
rect 17059 19245 17075 19279
rect 16790 19217 16824 19233
rect 16790 18833 16824 18849
rect 17118 19217 17152 19233
rect 17118 18833 17152 18849
rect 16867 18787 16883 18821
rect 17059 18787 17075 18821
rect 16672 18728 16748 18769
rect 17200 18769 17220 19297
rect 17254 18769 17330 19297
rect 17200 18728 17330 18769
rect 16672 18707 17330 18728
rect 16672 18673 16784 18707
rect 17158 18673 17330 18707
rect 16672 18643 17330 18673
rect 16672 18639 16748 18643
rect 16666 18128 16734 18129
rect 16850 18128 17330 18643
rect 16666 18103 17330 18128
rect 16666 18069 16784 18103
rect 17158 18069 17330 18103
rect 16666 18050 17330 18069
rect 16666 18007 16734 18050
rect 16666 17479 16688 18007
rect 16722 17479 16734 18007
rect 17200 18007 17330 18050
rect 16867 17955 16883 17989
rect 17059 17955 17075 17989
rect 16790 17927 16824 17943
rect 16790 17543 16824 17559
rect 17118 17927 17152 17943
rect 17118 17543 17152 17559
rect 16867 17497 16883 17531
rect 17059 17497 17075 17531
rect 16666 17438 16734 17479
rect 17200 17479 17220 18007
rect 17254 17490 17330 18007
rect 17469 17490 17624 22485
rect 22057 21625 22066 22815
rect 22404 22864 23955 22882
rect 22404 22830 22576 22864
rect 23832 22830 23955 22864
rect 22404 22815 23955 22830
rect 22404 22768 22540 22815
rect 22404 21982 22480 22768
rect 22514 21982 22540 22768
rect 23894 22768 23955 22815
rect 22650 22716 22666 22750
rect 23742 22716 23758 22750
rect 22582 22688 22616 22704
rect 22582 22404 22616 22420
rect 23792 22688 23826 22704
rect 23792 22404 23826 22420
rect 22650 22358 22666 22392
rect 23742 22358 23758 22392
rect 22582 22330 22616 22346
rect 22582 22046 22616 22062
rect 23792 22330 23826 22346
rect 23792 22046 23826 22062
rect 22650 22000 22666 22034
rect 23742 22000 23758 22034
rect 22404 21945 22540 21982
rect 23928 21982 23955 22768
rect 23894 21945 23955 21982
rect 22404 21920 23955 21945
rect 22404 21886 22576 21920
rect 23832 21886 23955 21920
rect 22404 21866 23955 21886
rect 24166 22878 24793 22882
rect 26051 22912 26057 23050
rect 26091 22912 26122 23050
rect 26051 22878 26122 22912
rect 24166 22850 26122 22878
rect 24166 22816 24855 22850
rect 25995 22816 26122 22850
rect 24166 22815 26122 22816
rect 22293 21625 23955 21627
rect 22057 21616 23955 21625
rect 24166 21616 24210 22815
rect 24283 22814 26122 22815
rect 22057 21565 24210 21616
rect 17254 17479 17624 17490
rect 17200 17438 17624 17479
rect 16666 17417 17624 17438
rect 16666 17383 16784 17417
rect 17158 17383 17624 17417
rect 16666 17362 17624 17383
rect 16668 17360 17624 17362
rect 15927 17060 16598 17074
rect 15106 17048 16598 17060
rect 15106 17014 15898 17048
rect 16480 17014 16598 17048
rect 17192 17029 17624 17360
rect 17192 17028 17429 17029
rect 17192 17017 17251 17028
rect 15106 16967 16598 17014
rect 16697 16968 16780 17017
rect 17159 16968 17251 17017
rect 15106 16962 15719 16967
rect 15106 16392 15242 16962
rect 16697 16906 16745 16968
rect 17192 16941 17251 16968
rect 16867 16867 16883 16901
rect 17059 16867 17075 16901
rect 17192 16899 17216 16941
rect 16790 16839 16824 16855
rect 16790 16655 16824 16671
rect 17118 16839 17152 16855
rect 17118 16655 17152 16671
rect 15106 16359 16524 16392
rect 15106 16325 15294 16359
rect 15328 16325 15384 16359
rect 15418 16325 15474 16359
rect 15508 16325 15564 16359
rect 15598 16325 15654 16359
rect 15688 16325 15744 16359
rect 15778 16325 15834 16359
rect 15868 16325 15924 16359
rect 15958 16325 16014 16359
rect 16048 16325 16104 16359
rect 16138 16325 16194 16359
rect 16228 16325 16284 16359
rect 16318 16325 16374 16359
rect 16408 16325 16524 16359
rect 15106 16316 16524 16325
rect 15106 16258 15334 16316
rect 15106 16224 15271 16258
rect 15305 16224 15334 16258
rect 15106 16208 15334 16224
rect 16377 16258 16524 16316
rect 16377 16224 16458 16258
rect 16492 16224 16524 16258
rect 16377 16208 16524 16224
rect 15106 16176 15494 16208
rect 15528 16176 15584 16208
rect 15618 16176 15674 16208
rect 15708 16176 15764 16208
rect 15798 16176 15854 16208
rect 15888 16176 15944 16208
rect 15978 16176 16034 16208
rect 16068 16176 16124 16208
rect 16158 16176 16214 16208
rect 16248 16176 16524 16208
rect 15106 16168 16524 16176
rect 15106 16134 15271 16168
rect 15305 16157 16458 16168
rect 15305 16152 15471 16157
rect 15305 16134 15418 16152
rect 15106 16118 15418 16134
rect 15452 16118 15471 16152
rect 15106 16078 15471 16118
rect 16289 16134 16458 16157
rect 16492 16134 16524 16168
rect 16289 16118 16524 16134
rect 15106 16044 15271 16078
rect 15305 16062 15471 16078
rect 15305 16044 15418 16062
rect 15106 16028 15418 16044
rect 15452 16028 15471 16062
rect 15106 15988 15471 16028
rect 15106 15954 15271 15988
rect 15305 15972 15471 15988
rect 15305 15954 15418 15972
rect 15106 15938 15418 15954
rect 15452 15938 15471 15972
rect 15106 15898 15471 15938
rect 15106 15864 15271 15898
rect 15305 15882 15471 15898
rect 15305 15864 15418 15882
rect 15106 15848 15418 15864
rect 15452 15848 15471 15882
rect 15106 15834 15471 15848
rect 15106 15315 15155 15834
rect 15019 15307 15155 15315
rect 15251 15808 15471 15834
rect 15251 15774 15271 15808
rect 15305 15792 15471 15808
rect 15305 15774 15418 15792
rect 15251 15758 15418 15774
rect 15452 15758 15471 15792
rect 15251 15718 15471 15758
rect 15251 15684 15271 15718
rect 15305 15702 15471 15718
rect 15305 15684 15418 15702
rect 15251 15668 15418 15684
rect 15452 15668 15471 15702
rect 15251 15628 15471 15668
rect 15251 15594 15271 15628
rect 15305 15612 15471 15628
rect 15305 15594 15418 15612
rect 15251 15578 15418 15594
rect 15452 15578 15471 15612
rect 15251 15538 15471 15578
rect 15251 15504 15271 15538
rect 15305 15522 15471 15538
rect 15305 15504 15418 15522
rect 15251 15488 15418 15504
rect 15452 15488 15471 15522
rect 15251 15448 15471 15488
rect 15251 15414 15271 15448
rect 15305 15432 15471 15448
rect 15305 15414 15418 15432
rect 15251 15398 15418 15414
rect 15452 15398 15471 15432
rect 15533 16036 16227 16095
rect 15533 16002 15592 16036
rect 15626 16008 15682 16036
rect 15654 16002 15682 16008
rect 15716 16008 15772 16036
rect 15716 16002 15720 16008
rect 15533 15974 15620 16002
rect 15654 15974 15720 16002
rect 15754 16002 15772 16008
rect 15806 16008 15862 16036
rect 15806 16002 15820 16008
rect 15754 15974 15820 16002
rect 15854 16002 15862 16008
rect 15896 16008 15952 16036
rect 15986 16008 16042 16036
rect 16076 16008 16132 16036
rect 15896 16002 15920 16008
rect 15986 16002 16020 16008
rect 16076 16002 16120 16008
rect 16166 16002 16227 16036
rect 15854 15974 15920 16002
rect 15954 15974 16020 16002
rect 16054 15974 16120 16002
rect 16154 15974 16227 16002
rect 15533 15946 16227 15974
rect 15533 15912 15592 15946
rect 15626 15912 15682 15946
rect 15716 15912 15772 15946
rect 15806 15912 15862 15946
rect 15896 15912 15952 15946
rect 15986 15912 16042 15946
rect 16076 15912 16132 15946
rect 16166 15912 16227 15946
rect 15533 15908 16227 15912
rect 15533 15874 15620 15908
rect 15654 15874 15720 15908
rect 15754 15874 15820 15908
rect 15854 15874 15920 15908
rect 15954 15874 16020 15908
rect 16054 15874 16120 15908
rect 16154 15874 16227 15908
rect 15533 15856 16227 15874
rect 15533 15822 15592 15856
rect 15626 15822 15682 15856
rect 15716 15822 15772 15856
rect 15806 15822 15862 15856
rect 15896 15822 15952 15856
rect 15986 15822 16042 15856
rect 16076 15822 16132 15856
rect 16166 15822 16227 15856
rect 15533 15808 16227 15822
rect 15533 15774 15620 15808
rect 15654 15774 15720 15808
rect 15754 15774 15820 15808
rect 15854 15774 15920 15808
rect 15954 15774 16020 15808
rect 16054 15774 16120 15808
rect 16154 15774 16227 15808
rect 15533 15766 16227 15774
rect 15533 15732 15592 15766
rect 15626 15732 15682 15766
rect 15716 15732 15772 15766
rect 15806 15732 15862 15766
rect 15896 15732 15952 15766
rect 15986 15732 16042 15766
rect 16076 15732 16132 15766
rect 16166 15732 16227 15766
rect 15533 15708 16227 15732
rect 15533 15676 15620 15708
rect 15654 15676 15720 15708
rect 15533 15642 15592 15676
rect 15654 15674 15682 15676
rect 15626 15642 15682 15674
rect 15716 15674 15720 15676
rect 15754 15676 15820 15708
rect 15754 15674 15772 15676
rect 15716 15642 15772 15674
rect 15806 15674 15820 15676
rect 15854 15676 15920 15708
rect 15954 15676 16020 15708
rect 16054 15676 16120 15708
rect 16154 15676 16227 15708
rect 15854 15674 15862 15676
rect 15806 15642 15862 15674
rect 15896 15674 15920 15676
rect 15986 15674 16020 15676
rect 16076 15674 16120 15676
rect 15896 15642 15952 15674
rect 15986 15642 16042 15674
rect 16076 15642 16132 15674
rect 16166 15642 16227 15676
rect 15533 15608 16227 15642
rect 15533 15586 15620 15608
rect 15654 15586 15720 15608
rect 15533 15552 15592 15586
rect 15654 15574 15682 15586
rect 15626 15552 15682 15574
rect 15716 15574 15720 15586
rect 15754 15586 15820 15608
rect 15754 15574 15772 15586
rect 15716 15552 15772 15574
rect 15806 15574 15820 15586
rect 15854 15586 15920 15608
rect 15954 15586 16020 15608
rect 16054 15586 16120 15608
rect 16154 15586 16227 15608
rect 15854 15574 15862 15586
rect 15806 15552 15862 15574
rect 15896 15574 15920 15586
rect 15986 15574 16020 15586
rect 16076 15574 16120 15586
rect 15896 15552 15952 15574
rect 15986 15552 16042 15574
rect 16076 15552 16132 15574
rect 16166 15552 16227 15586
rect 15533 15508 16227 15552
rect 15533 15496 15620 15508
rect 15654 15496 15720 15508
rect 15533 15462 15592 15496
rect 15654 15474 15682 15496
rect 15626 15462 15682 15474
rect 15716 15474 15720 15496
rect 15754 15496 15820 15508
rect 15754 15474 15772 15496
rect 15716 15462 15772 15474
rect 15806 15474 15820 15496
rect 15854 15496 15920 15508
rect 15954 15496 16020 15508
rect 16054 15496 16120 15508
rect 16154 15496 16227 15508
rect 15854 15474 15862 15496
rect 15806 15462 15862 15474
rect 15896 15474 15920 15496
rect 15986 15474 16020 15496
rect 16076 15474 16120 15496
rect 15896 15462 15952 15474
rect 15986 15462 16042 15474
rect 16076 15462 16132 15474
rect 16166 15462 16227 15496
rect 15533 15401 16227 15462
rect 16289 16084 16308 16118
rect 16342 16084 16524 16118
rect 16289 16083 16524 16084
rect 16289 16028 16344 16083
rect 16289 15994 16308 16028
rect 16342 15994 16344 16028
rect 16289 15938 16344 15994
rect 16289 15904 16308 15938
rect 16342 15904 16344 15938
rect 16289 15848 16344 15904
rect 16289 15814 16308 15848
rect 16342 15814 16344 15848
rect 16289 15758 16344 15814
rect 16289 15724 16308 15758
rect 16342 15724 16344 15758
rect 16289 15668 16344 15724
rect 16289 15634 16308 15668
rect 16342 15634 16344 15668
rect 16289 15578 16344 15634
rect 16289 15544 16308 15578
rect 16342 15544 16344 15578
rect 16289 15488 16344 15544
rect 16289 15454 16308 15488
rect 16342 15454 16344 15488
rect 15251 15358 15471 15398
rect 15251 15324 15271 15358
rect 15305 15339 15471 15358
rect 16289 15398 16344 15454
rect 16289 15364 16308 15398
rect 16342 15364 16344 15398
rect 16289 15339 16344 15364
rect 15305 15324 16344 15339
rect 15251 15320 16344 15324
rect 15251 15307 15475 15320
rect 15019 15286 15475 15307
rect 15509 15286 15565 15320
rect 15599 15286 15655 15320
rect 15689 15286 15745 15320
rect 15779 15286 15835 15320
rect 15869 15286 15925 15320
rect 15959 15286 16015 15320
rect 16049 15286 16105 15320
rect 16139 15286 16195 15320
rect 16229 15286 16344 15320
rect 15019 15281 16344 15286
rect 15019 15268 15767 15281
rect 15019 15234 15271 15268
rect 15305 15234 15767 15268
rect 15019 15198 15767 15234
rect 12227 15179 15767 15198
rect 12227 15172 12309 15179
rect 12461 15172 13299 15179
rect 13447 15172 15767 15179
rect 16246 15258 16344 15281
rect 16246 15234 16458 15258
rect 16492 15234 16524 16083
rect 16246 15172 16524 15234
rect 12227 15138 12250 15172
rect 14959 15138 15294 15172
rect 15328 15138 15384 15172
rect 15418 15138 15474 15172
rect 15508 15138 15564 15172
rect 15598 15138 15654 15172
rect 15688 15138 15744 15172
rect 16246 15161 16284 15172
rect 15778 15138 15834 15161
rect 15868 15138 15924 15161
rect 15958 15138 16014 15161
rect 16048 15138 16104 15161
rect 16138 15138 16194 15161
rect 16228 15138 16284 15161
rect 16318 15138 16374 15172
rect 16408 15138 16524 15172
rect 12227 15125 12309 15138
rect 12461 15125 13299 15138
rect 13447 15125 16524 15138
rect 12227 15122 16524 15125
rect 11975 15106 16524 15122
rect 11975 15019 12336 15106
rect 15150 15105 16524 15106
rect 15236 15104 16524 15105
rect 16697 16372 16745 16629
rect 16867 16609 16883 16643
rect 17059 16609 17075 16643
rect 16790 16581 16824 16597
rect 16790 16397 16824 16413
rect 17118 16581 17152 16597
rect 17118 16397 17152 16413
rect 16867 16351 16883 16385
rect 17059 16351 17075 16385
rect 17192 16273 17195 16899
rect 16867 16142 16883 16176
rect 16959 16142 16975 16176
rect 16790 16114 16824 16130
rect 16790 15730 16824 15746
rect 17018 16114 17052 16130
rect 17018 15730 17052 15746
rect 16867 15684 16883 15718
rect 16959 15684 16975 15718
rect 16790 15656 16824 15672
rect 16790 15272 16824 15288
rect 17018 15656 17052 15672
rect 17018 15272 17052 15288
rect 17189 15285 17195 16273
rect 17351 16042 17429 17028
rect 16697 15128 16745 15264
rect 16867 15226 16883 15260
rect 16959 15226 16975 15260
rect 17190 15239 17195 15285
rect 17189 15224 17195 15239
rect 17189 15128 17218 15224
rect 16697 15076 16864 15128
rect 17100 15076 17218 15128
rect 17189 15049 17218 15076
rect 17350 15050 17429 16042
rect 17577 16925 17624 17029
rect 17577 15050 17623 16925
rect 17350 15049 17623 15050
rect 17189 14999 17623 15049
rect 17726 11104 25902 11140
rect 17726 11015 17910 11104
rect 25708 11015 25902 11104
rect 17726 10959 25902 11015
rect 17726 10925 17978 10959
rect 25666 10925 25902 10959
rect 17726 10899 25902 10925
rect 2610 10423 2971 10510
rect 7824 10480 8258 10530
rect 7824 10453 7853 10480
rect 5871 10424 7159 10425
rect 5785 10423 7159 10424
rect 2610 10407 7159 10423
rect 2610 3829 2688 10407
rect 2862 10404 7159 10407
rect 2862 10391 2944 10404
rect 3096 10391 3934 10404
rect 4082 10391 7159 10404
rect 2862 10357 2885 10391
rect 5594 10357 5929 10391
rect 5963 10357 6019 10391
rect 6053 10357 6109 10391
rect 6143 10357 6199 10391
rect 6233 10357 6289 10391
rect 6323 10357 6379 10391
rect 6413 10368 6469 10391
rect 6503 10368 6559 10391
rect 6593 10368 6649 10391
rect 6683 10368 6739 10391
rect 6773 10368 6829 10391
rect 6863 10368 6919 10391
rect 6881 10357 6919 10368
rect 6953 10357 7009 10391
rect 7043 10357 7159 10391
rect 2862 10350 2944 10357
rect 3096 10350 3934 10357
rect 4082 10350 6402 10357
rect 2862 10331 6402 10350
rect 2862 3908 2971 10331
rect 3097 10151 3113 10185
rect 3889 10151 3905 10185
rect 4578 10151 4594 10185
rect 5370 10151 5386 10185
rect 5584 10171 5620 10331
rect 5654 10295 6402 10331
rect 5654 10261 5906 10295
rect 5940 10261 6402 10295
rect 5654 10248 6402 10261
rect 6881 10295 7159 10357
rect 6881 10271 7093 10295
rect 6881 10248 6979 10271
rect 5654 10243 6979 10248
rect 5654 10222 6110 10243
rect 5654 10214 5790 10222
rect 3029 10123 3063 10139
rect 3029 9939 3063 9955
rect 3939 10123 3973 10139
rect 3939 9939 3973 9955
rect 4510 10123 4544 10139
rect 4510 9939 4544 9955
rect 5420 10123 5454 10139
rect 5420 9939 5454 9955
rect 3097 9893 3113 9927
rect 3889 9893 3905 9927
rect 4578 9893 4594 9927
rect 5370 9893 5386 9927
rect 3029 9865 3063 9881
rect 3029 9681 3063 9697
rect 3939 9865 3973 9881
rect 3939 9681 3973 9697
rect 4510 9865 4544 9881
rect 4510 9681 4544 9697
rect 5420 9865 5454 9881
rect 5420 9681 5454 9697
rect 3097 9635 3113 9669
rect 3889 9635 3905 9669
rect 4578 9635 4594 9669
rect 5370 9635 5386 9669
rect 3029 9607 3063 9623
rect 3029 9423 3063 9439
rect 3939 9607 3973 9623
rect 3939 9423 3973 9439
rect 4510 9607 4544 9623
rect 4510 9423 4544 9439
rect 5420 9607 5454 9623
rect 5420 9423 5454 9439
rect 3097 9377 3113 9411
rect 3889 9377 3905 9411
rect 4578 9377 4594 9411
rect 5370 9377 5386 9411
rect 3029 9349 3063 9365
rect 3029 9165 3063 9181
rect 3939 9349 3973 9365
rect 3939 9165 3973 9181
rect 4510 9349 4544 9365
rect 4510 9165 4544 9181
rect 5420 9349 5454 9365
rect 5420 9165 5454 9181
rect 3097 9119 3113 9153
rect 3889 9119 3905 9153
rect 4578 9119 4594 9153
rect 5370 9119 5386 9153
rect 3029 9091 3063 9107
rect 3029 8907 3063 8923
rect 3939 9091 3973 9107
rect 3939 8907 3973 8923
rect 4510 9091 4544 9107
rect 4510 8907 4544 8923
rect 5420 9091 5454 9107
rect 5420 8907 5454 8923
rect 3097 8861 3113 8895
rect 3889 8861 3905 8895
rect 4578 8861 4594 8895
rect 5370 8861 5386 8895
rect 3029 8833 3063 8849
rect 3029 8649 3063 8665
rect 3939 8833 3973 8849
rect 3939 8649 3973 8665
rect 4510 8833 4544 8849
rect 4510 8649 4544 8665
rect 5420 8833 5454 8849
rect 5420 8649 5454 8665
rect 3097 8603 3113 8637
rect 3889 8603 3905 8637
rect 4578 8603 4594 8637
rect 5370 8603 5386 8637
rect 3029 8575 3063 8591
rect 3029 8391 3063 8407
rect 3939 8575 3973 8591
rect 3939 8391 3973 8407
rect 4510 8575 4544 8591
rect 4510 8391 4544 8407
rect 5420 8575 5454 8591
rect 5420 8391 5454 8407
rect 3097 8345 3113 8379
rect 3889 8345 3905 8379
rect 4578 8345 4594 8379
rect 5370 8345 5386 8379
rect 3029 8317 3063 8333
rect 3029 8133 3063 8149
rect 3939 8317 3973 8333
rect 3939 8133 3973 8149
rect 4510 8317 4544 8333
rect 4510 8133 4544 8149
rect 5420 8317 5454 8333
rect 5420 8133 5454 8149
rect 3097 8087 3113 8121
rect 3889 8087 3905 8121
rect 4578 8087 4594 8121
rect 5370 8087 5386 8121
rect 3029 8059 3063 8075
rect 3029 7875 3063 7891
rect 3939 8059 3973 8075
rect 3939 7875 3973 7891
rect 4510 8059 4544 8075
rect 4510 7875 4544 7891
rect 5420 8059 5454 8075
rect 5420 7875 5454 7891
rect 3097 7829 3113 7863
rect 3889 7829 3905 7863
rect 4578 7829 4594 7863
rect 5370 7829 5386 7863
rect 3029 7801 3063 7817
rect 3029 7617 3063 7633
rect 3939 7801 3973 7817
rect 3939 7617 3973 7633
rect 4510 7801 4544 7817
rect 4510 7617 4544 7633
rect 5420 7801 5454 7817
rect 5420 7617 5454 7633
rect 3097 7571 3113 7605
rect 3889 7571 3905 7605
rect 4578 7571 4594 7605
rect 5370 7571 5386 7605
rect 3029 7543 3063 7559
rect 3029 7359 3063 7375
rect 3939 7543 3973 7559
rect 3939 7359 3973 7375
rect 4510 7543 4544 7559
rect 4510 7359 4544 7375
rect 5420 7543 5454 7559
rect 5420 7359 5454 7375
rect 3097 7313 3113 7347
rect 3889 7313 3905 7347
rect 4578 7313 4594 7347
rect 5370 7313 5386 7347
rect 3029 7285 3063 7301
rect 3029 7101 3063 7117
rect 3939 7285 3973 7301
rect 3939 7101 3973 7117
rect 4510 7285 4544 7301
rect 4510 7101 4544 7117
rect 5420 7285 5454 7301
rect 5420 7101 5454 7117
rect 3097 7055 3113 7089
rect 3889 7055 3905 7089
rect 4578 7055 4594 7089
rect 5370 7055 5386 7089
rect 3029 7027 3063 7043
rect 3029 6843 3063 6859
rect 3939 7027 3973 7043
rect 3939 6843 3973 6859
rect 4510 7027 4544 7043
rect 4510 6843 4544 6859
rect 5420 7027 5454 7043
rect 5420 6843 5454 6859
rect 3097 6797 3113 6831
rect 3889 6797 3905 6831
rect 4578 6797 4594 6831
rect 5370 6797 5386 6831
rect 3029 6769 3063 6785
rect 3029 6585 3063 6601
rect 3939 6769 3973 6785
rect 3939 6585 3973 6601
rect 4510 6769 4544 6785
rect 4510 6585 4544 6601
rect 5420 6769 5454 6785
rect 5420 6585 5454 6601
rect 3097 6539 3113 6573
rect 3889 6539 3905 6573
rect 4578 6539 4594 6573
rect 5370 6539 5386 6573
rect 3029 6511 3063 6527
rect 3029 6327 3063 6343
rect 3939 6511 3973 6527
rect 3939 6327 3973 6343
rect 4510 6511 4544 6527
rect 4510 6327 4544 6343
rect 5420 6511 5454 6527
rect 5420 6327 5454 6343
rect 3097 6281 3113 6315
rect 3889 6281 3905 6315
rect 4578 6281 4594 6315
rect 5370 6281 5386 6315
rect 3029 6253 3063 6269
rect 3029 6069 3063 6085
rect 3939 6253 3973 6269
rect 3939 6069 3973 6085
rect 4510 6253 4544 6269
rect 4510 6069 4544 6085
rect 5420 6253 5454 6269
rect 5420 6069 5454 6085
rect 3097 6023 3113 6057
rect 3889 6023 3905 6057
rect 4578 6023 4594 6057
rect 5370 6023 5386 6057
rect 3029 5995 3063 6011
rect 3029 5811 3063 5827
rect 3939 5995 3973 6011
rect 3939 5811 3973 5827
rect 4510 5995 4544 6011
rect 4510 5811 4544 5827
rect 5420 5995 5454 6011
rect 5420 5811 5454 5827
rect 3097 5765 3113 5799
rect 3889 5765 3905 5799
rect 4578 5765 4594 5799
rect 5370 5765 5386 5799
rect 3029 5737 3063 5753
rect 3029 5553 3063 5569
rect 3939 5737 3973 5753
rect 3939 5553 3973 5569
rect 4510 5737 4544 5753
rect 4510 5553 4544 5569
rect 5420 5737 5454 5753
rect 5420 5553 5454 5569
rect 3097 5507 3113 5541
rect 3889 5507 3905 5541
rect 4578 5507 4594 5541
rect 5370 5507 5386 5541
rect 3029 5479 3063 5495
rect 3029 5295 3063 5311
rect 3939 5479 3973 5495
rect 3939 5295 3973 5311
rect 4510 5479 4544 5495
rect 4510 5295 4544 5311
rect 5420 5479 5454 5495
rect 5420 5295 5454 5311
rect 3097 5249 3113 5283
rect 3889 5249 3905 5283
rect 4578 5249 4594 5283
rect 5370 5249 5386 5283
rect 3029 5221 3063 5237
rect 3029 5037 3063 5053
rect 3939 5221 3973 5237
rect 3939 5037 3973 5053
rect 4510 5221 4544 5237
rect 4510 5037 4544 5053
rect 5420 5221 5454 5237
rect 5420 5037 5454 5053
rect 3097 4991 3113 5025
rect 3889 4991 3905 5025
rect 4578 4991 4594 5025
rect 5370 4991 5386 5025
rect 3029 4963 3063 4979
rect 3029 4779 3063 4795
rect 3939 4963 3973 4979
rect 3939 4779 3973 4795
rect 4510 4963 4544 4979
rect 4510 4779 4544 4795
rect 5420 4963 5454 4979
rect 5420 4779 5454 4795
rect 3097 4733 3113 4767
rect 3889 4733 3905 4767
rect 4578 4733 4594 4767
rect 5370 4733 5386 4767
rect 3029 4705 3063 4721
rect 3029 4521 3063 4537
rect 3939 4705 3973 4721
rect 3939 4521 3973 4537
rect 4510 4705 4544 4721
rect 4510 4521 4544 4537
rect 5420 4705 5454 4721
rect 5420 4521 5454 4537
rect 3097 4475 3113 4509
rect 3889 4475 3905 4509
rect 4578 4475 4594 4509
rect 5370 4475 5386 4509
rect 3029 4447 3063 4463
rect 3029 4263 3063 4279
rect 3939 4447 3973 4463
rect 3939 4263 3973 4279
rect 4510 4447 4544 4463
rect 4510 4263 4544 4279
rect 5420 4447 5454 4463
rect 5420 4263 5454 4279
rect 3097 4217 3113 4251
rect 3889 4217 3905 4251
rect 4578 4217 4594 4251
rect 5370 4217 5386 4251
rect 3029 4189 3063 4205
rect 3029 4005 3063 4021
rect 3939 4189 3973 4205
rect 3939 4005 3973 4021
rect 4510 4189 4544 4205
rect 4510 4005 4544 4021
rect 5420 4189 5454 4205
rect 5420 4005 5454 4021
rect 3097 3959 3113 3993
rect 3889 3959 3905 3993
rect 4578 3959 4594 3993
rect 5370 3959 5386 3993
rect 5577 3908 5620 10171
rect 2862 3875 5620 3908
rect 5741 9695 5790 10214
rect 5886 10209 6110 10222
rect 6144 10209 6200 10243
rect 6234 10209 6290 10243
rect 6324 10209 6380 10243
rect 6414 10209 6470 10243
rect 6504 10209 6560 10243
rect 6594 10209 6650 10243
rect 6684 10209 6740 10243
rect 6774 10209 6830 10243
rect 6864 10209 6979 10243
rect 5886 10205 6979 10209
rect 5886 10171 5906 10205
rect 5940 10190 6979 10205
rect 5940 10171 6106 10190
rect 5886 10131 6106 10171
rect 5886 10115 6053 10131
rect 5886 10081 5906 10115
rect 5940 10097 6053 10115
rect 6087 10097 6106 10131
rect 6924 10165 6979 10190
rect 6924 10131 6943 10165
rect 6977 10131 6979 10165
rect 5940 10081 6106 10097
rect 5886 10041 6106 10081
rect 5886 10025 6053 10041
rect 5886 9991 5906 10025
rect 5940 10007 6053 10025
rect 6087 10007 6106 10041
rect 5940 9991 6106 10007
rect 5886 9951 6106 9991
rect 5886 9935 6053 9951
rect 5886 9901 5906 9935
rect 5940 9917 6053 9935
rect 6087 9917 6106 9951
rect 5940 9901 6106 9917
rect 5886 9861 6106 9901
rect 5886 9845 6053 9861
rect 5886 9811 5906 9845
rect 5940 9827 6053 9845
rect 6087 9827 6106 9861
rect 5940 9811 6106 9827
rect 5886 9771 6106 9811
rect 5886 9755 6053 9771
rect 5886 9721 5906 9755
rect 5940 9737 6053 9755
rect 6087 9737 6106 9771
rect 5940 9721 6106 9737
rect 5886 9695 6106 9721
rect 5741 9681 6106 9695
rect 5741 9665 6053 9681
rect 5741 9631 5906 9665
rect 5940 9647 6053 9665
rect 6087 9647 6106 9681
rect 5940 9631 6106 9647
rect 5741 9591 6106 9631
rect 5741 9575 6053 9591
rect 5741 9541 5906 9575
rect 5940 9557 6053 9575
rect 6087 9557 6106 9591
rect 5940 9541 6106 9557
rect 5741 9501 6106 9541
rect 5741 9485 6053 9501
rect 5741 9451 5906 9485
rect 5940 9467 6053 9485
rect 6087 9467 6106 9501
rect 5940 9451 6106 9467
rect 5741 9411 6106 9451
rect 6168 10067 6862 10128
rect 6168 10033 6227 10067
rect 6261 10055 6317 10067
rect 6289 10033 6317 10055
rect 6351 10055 6407 10067
rect 6351 10033 6355 10055
rect 6168 10021 6255 10033
rect 6289 10021 6355 10033
rect 6389 10033 6407 10055
rect 6441 10055 6497 10067
rect 6441 10033 6455 10055
rect 6389 10021 6455 10033
rect 6489 10033 6497 10055
rect 6531 10055 6587 10067
rect 6621 10055 6677 10067
rect 6711 10055 6767 10067
rect 6531 10033 6555 10055
rect 6621 10033 6655 10055
rect 6711 10033 6755 10055
rect 6801 10033 6862 10067
rect 6489 10021 6555 10033
rect 6589 10021 6655 10033
rect 6689 10021 6755 10033
rect 6789 10021 6862 10033
rect 6168 9977 6862 10021
rect 6168 9943 6227 9977
rect 6261 9955 6317 9977
rect 6289 9943 6317 9955
rect 6351 9955 6407 9977
rect 6351 9943 6355 9955
rect 6168 9921 6255 9943
rect 6289 9921 6355 9943
rect 6389 9943 6407 9955
rect 6441 9955 6497 9977
rect 6441 9943 6455 9955
rect 6389 9921 6455 9943
rect 6489 9943 6497 9955
rect 6531 9955 6587 9977
rect 6621 9955 6677 9977
rect 6711 9955 6767 9977
rect 6531 9943 6555 9955
rect 6621 9943 6655 9955
rect 6711 9943 6755 9955
rect 6801 9943 6862 9977
rect 6489 9921 6555 9943
rect 6589 9921 6655 9943
rect 6689 9921 6755 9943
rect 6789 9921 6862 9943
rect 6168 9887 6862 9921
rect 6168 9853 6227 9887
rect 6261 9855 6317 9887
rect 6289 9853 6317 9855
rect 6351 9855 6407 9887
rect 6351 9853 6355 9855
rect 6168 9821 6255 9853
rect 6289 9821 6355 9853
rect 6389 9853 6407 9855
rect 6441 9855 6497 9887
rect 6441 9853 6455 9855
rect 6389 9821 6455 9853
rect 6489 9853 6497 9855
rect 6531 9855 6587 9887
rect 6621 9855 6677 9887
rect 6711 9855 6767 9887
rect 6531 9853 6555 9855
rect 6621 9853 6655 9855
rect 6711 9853 6755 9855
rect 6801 9853 6862 9887
rect 6489 9821 6555 9853
rect 6589 9821 6655 9853
rect 6689 9821 6755 9853
rect 6789 9821 6862 9853
rect 6168 9797 6862 9821
rect 6168 9763 6227 9797
rect 6261 9763 6317 9797
rect 6351 9763 6407 9797
rect 6441 9763 6497 9797
rect 6531 9763 6587 9797
rect 6621 9763 6677 9797
rect 6711 9763 6767 9797
rect 6801 9763 6862 9797
rect 6168 9755 6862 9763
rect 6168 9721 6255 9755
rect 6289 9721 6355 9755
rect 6389 9721 6455 9755
rect 6489 9721 6555 9755
rect 6589 9721 6655 9755
rect 6689 9721 6755 9755
rect 6789 9721 6862 9755
rect 6168 9707 6862 9721
rect 6168 9673 6227 9707
rect 6261 9673 6317 9707
rect 6351 9673 6407 9707
rect 6441 9673 6497 9707
rect 6531 9673 6587 9707
rect 6621 9673 6677 9707
rect 6711 9673 6767 9707
rect 6801 9673 6862 9707
rect 6168 9655 6862 9673
rect 6168 9621 6255 9655
rect 6289 9621 6355 9655
rect 6389 9621 6455 9655
rect 6489 9621 6555 9655
rect 6589 9621 6655 9655
rect 6689 9621 6755 9655
rect 6789 9621 6862 9655
rect 6168 9617 6862 9621
rect 6168 9583 6227 9617
rect 6261 9583 6317 9617
rect 6351 9583 6407 9617
rect 6441 9583 6497 9617
rect 6531 9583 6587 9617
rect 6621 9583 6677 9617
rect 6711 9583 6767 9617
rect 6801 9583 6862 9617
rect 6168 9555 6862 9583
rect 6168 9527 6255 9555
rect 6289 9527 6355 9555
rect 6168 9493 6227 9527
rect 6289 9521 6317 9527
rect 6261 9493 6317 9521
rect 6351 9521 6355 9527
rect 6389 9527 6455 9555
rect 6389 9521 6407 9527
rect 6351 9493 6407 9521
rect 6441 9521 6455 9527
rect 6489 9527 6555 9555
rect 6589 9527 6655 9555
rect 6689 9527 6755 9555
rect 6789 9527 6862 9555
rect 6489 9521 6497 9527
rect 6441 9493 6497 9521
rect 6531 9521 6555 9527
rect 6621 9521 6655 9527
rect 6711 9521 6755 9527
rect 6531 9493 6587 9521
rect 6621 9493 6677 9521
rect 6711 9493 6767 9521
rect 6801 9493 6862 9527
rect 6168 9434 6862 9493
rect 6924 10075 6979 10131
rect 6924 10041 6943 10075
rect 6977 10041 6979 10075
rect 6924 9985 6979 10041
rect 6924 9951 6943 9985
rect 6977 9951 6979 9985
rect 6924 9895 6979 9951
rect 6924 9861 6943 9895
rect 6977 9861 6979 9895
rect 6924 9805 6979 9861
rect 6924 9771 6943 9805
rect 6977 9771 6979 9805
rect 6924 9715 6979 9771
rect 6924 9681 6943 9715
rect 6977 9681 6979 9715
rect 6924 9625 6979 9681
rect 6924 9591 6943 9625
rect 6977 9591 6979 9625
rect 6924 9535 6979 9591
rect 6924 9501 6943 9535
rect 6977 9501 6979 9535
rect 6924 9446 6979 9501
rect 7127 9446 7159 10295
rect 6924 9445 7159 9446
rect 5741 9395 6053 9411
rect 5741 9361 5906 9395
rect 5940 9377 6053 9395
rect 6087 9377 6106 9411
rect 5940 9372 6106 9377
rect 6924 9411 6943 9445
rect 6977 9411 7159 9445
rect 6924 9395 7159 9411
rect 6924 9372 7093 9395
rect 5940 9361 7093 9372
rect 7127 9361 7159 9395
rect 5741 9353 7159 9361
rect 5741 9321 6129 9353
rect 6163 9321 6219 9353
rect 6253 9321 6309 9353
rect 6343 9321 6399 9353
rect 6433 9321 6489 9353
rect 6523 9321 6579 9353
rect 6613 9321 6669 9353
rect 6703 9321 6759 9353
rect 6793 9321 6849 9353
rect 6883 9321 7159 9353
rect 5741 9305 5969 9321
rect 5741 9271 5906 9305
rect 5940 9271 5969 9305
rect 5741 9213 5969 9271
rect 7012 9305 7159 9321
rect 7012 9271 7093 9305
rect 7127 9271 7159 9305
rect 7012 9213 7159 9271
rect 5741 9204 7159 9213
rect 5741 9170 5929 9204
rect 5963 9170 6019 9204
rect 6053 9170 6109 9204
rect 6143 9170 6199 9204
rect 6233 9170 6289 9204
rect 6323 9170 6379 9204
rect 6413 9170 6469 9204
rect 6503 9170 6559 9204
rect 6593 9170 6649 9204
rect 6683 9170 6739 9204
rect 6773 9170 6829 9204
rect 6863 9170 6919 9204
rect 6953 9170 7009 9204
rect 7043 9170 7159 9204
rect 5741 9137 7159 9170
rect 7332 10401 7499 10453
rect 7735 10401 7853 10453
rect 7332 10265 7380 10401
rect 7824 10305 7853 10401
rect 7985 10479 8258 10480
rect 7502 10269 7518 10303
rect 7594 10269 7610 10303
rect 7824 10290 7830 10305
rect 7425 10241 7459 10257
rect 7425 9857 7459 9873
rect 7653 10241 7687 10257
rect 7825 10244 7830 10290
rect 7653 9857 7687 9873
rect 7502 9811 7518 9845
rect 7594 9811 7610 9845
rect 7425 9783 7459 9799
rect 7425 9399 7459 9415
rect 7653 9783 7687 9799
rect 7653 9399 7687 9415
rect 7502 9353 7518 9387
rect 7594 9353 7610 9387
rect 7824 9256 7830 10244
rect 7985 9487 8064 10479
rect 5741 8464 5877 9137
rect 7332 8900 7380 9157
rect 7502 9144 7518 9178
rect 7694 9144 7710 9178
rect 7425 9116 7459 9132
rect 7425 8932 7459 8948
rect 7753 9116 7787 9132
rect 7753 8932 7787 8948
rect 7502 8886 7518 8920
rect 7694 8886 7710 8920
rect 7425 8858 7459 8874
rect 7425 8674 7459 8690
rect 7753 8858 7787 8874
rect 7753 8674 7787 8690
rect 7502 8628 7518 8662
rect 7694 8628 7710 8662
rect 7827 8630 7830 9256
rect 7332 8561 7380 8623
rect 7827 8588 7851 8630
rect 7827 8561 7886 8588
rect 7332 8512 7415 8561
rect 7794 8512 7886 8561
rect 7827 8501 7886 8512
rect 7986 8501 8064 9487
rect 7827 8500 8064 8501
rect 8212 8500 8258 10479
rect 17726 9643 17918 10899
rect 17952 10802 25692 10899
rect 17952 9643 17980 10802
rect 18221 10713 18237 10747
rect 21805 10713 21821 10747
rect 21879 10713 21895 10747
rect 25463 10713 25479 10747
rect 18175 10654 18209 10670
rect 18175 10302 18209 10318
rect 21833 10654 21867 10670
rect 21833 10302 21867 10318
rect 25491 10654 25525 10670
rect 25491 10302 25525 10318
rect 18221 10225 18237 10259
rect 21805 10225 21821 10259
rect 21879 10225 21895 10259
rect 25463 10225 25479 10259
rect 18175 10166 18209 10182
rect 18175 9814 18209 9830
rect 21833 10166 21867 10182
rect 21833 9814 21867 9830
rect 25491 10166 25525 10182
rect 25491 9814 25525 9830
rect 18221 9737 18237 9771
rect 21805 9737 21821 9771
rect 21879 9737 21895 9771
rect 25463 9737 25479 9771
rect 17726 9633 17980 9643
rect 25726 10802 25902 10899
rect 25726 9643 25901 10802
rect 25692 9633 25901 9643
rect 17726 9617 25901 9633
rect 17726 9583 17978 9617
rect 25666 9583 25901 9617
rect 17726 9500 25901 9583
rect 7827 8477 8258 8500
rect 17727 8998 24876 9065
rect 17727 8964 19209 8998
rect 24510 8964 24876 8998
rect 17727 8938 24876 8964
rect 5741 8463 6352 8464
rect 5741 8416 7233 8463
rect 5741 8382 6533 8416
rect 7115 8382 7233 8416
rect 5741 8370 7233 8382
rect 2862 3873 5629 3875
rect 5741 3873 6371 8370
rect 6562 8356 7233 8370
rect 2862 3849 6371 3873
rect 2862 3829 2885 3849
rect 2610 3815 2885 3829
rect 5594 3815 6371 3849
rect 2610 3792 6371 3815
rect 6343 2963 6371 3792
rect 6562 8340 7141 8356
rect 6562 2964 6599 8340
rect 6715 8215 6731 8249
rect 6907 8215 6923 8249
rect 6647 8187 6681 8203
rect 6647 8003 6681 8019
rect 6957 8187 6991 8203
rect 6957 8003 6991 8019
rect 6715 7957 6731 7991
rect 6907 7957 6923 7991
rect 6647 7929 6681 7945
rect 6647 7745 6681 7761
rect 6957 7929 6991 7945
rect 6957 7745 6991 7761
rect 6715 7699 6731 7733
rect 6907 7699 6923 7733
rect 6647 7671 6681 7687
rect 6647 7487 6681 7503
rect 6957 7671 6991 7687
rect 6957 7487 6991 7503
rect 6715 7441 6731 7475
rect 6907 7441 6923 7475
rect 6647 7413 6681 7429
rect 6647 7229 6681 7245
rect 6957 7413 6991 7429
rect 6957 7229 6991 7245
rect 6715 7183 6731 7217
rect 6907 7183 6923 7217
rect 6647 7155 6681 7171
rect 6647 6971 6681 6987
rect 6957 7155 6991 7171
rect 6957 6971 6991 6987
rect 6715 6925 6731 6959
rect 6907 6925 6923 6959
rect 6647 6897 6681 6913
rect 6647 6713 6681 6729
rect 6957 6897 6991 6913
rect 6957 6713 6991 6729
rect 6715 6667 6731 6701
rect 6907 6667 6923 6701
rect 6647 6639 6681 6655
rect 6647 6455 6681 6471
rect 6957 6639 6991 6655
rect 6957 6455 6991 6471
rect 6715 6409 6731 6443
rect 6907 6409 6923 6443
rect 6647 6381 6681 6397
rect 6647 6197 6681 6213
rect 6957 6381 6991 6397
rect 6957 6197 6991 6213
rect 6715 6151 6731 6185
rect 6907 6151 6923 6185
rect 6647 6123 6681 6139
rect 6647 5939 6681 5955
rect 6957 6123 6991 6139
rect 6957 5939 6991 5955
rect 6715 5893 6731 5927
rect 6907 5893 6923 5927
rect 6647 5865 6681 5881
rect 6647 5681 6681 5697
rect 6957 5865 6991 5881
rect 6957 5681 6991 5697
rect 6715 5635 6731 5669
rect 6907 5635 6923 5669
rect 6647 5607 6681 5623
rect 6647 5423 6681 5439
rect 6957 5607 6991 5623
rect 6957 5423 6991 5439
rect 6715 5377 6731 5411
rect 6907 5377 6923 5411
rect 6647 5349 6681 5365
rect 6647 5165 6681 5181
rect 6957 5349 6991 5365
rect 6957 5165 6991 5181
rect 6715 5119 6731 5153
rect 6907 5119 6923 5153
rect 6647 5091 6681 5107
rect 6647 4907 6681 4923
rect 6957 5091 6991 5107
rect 6957 4907 6991 4923
rect 6715 4861 6731 4895
rect 6907 4861 6923 4895
rect 6647 4833 6681 4849
rect 6647 4649 6681 4665
rect 6957 4833 6991 4849
rect 6957 4649 6991 4665
rect 6715 4603 6731 4637
rect 6907 4603 6923 4637
rect 6647 4575 6681 4591
rect 6647 4391 6681 4407
rect 6957 4575 6991 4591
rect 6957 4391 6991 4407
rect 6715 4345 6731 4379
rect 6907 4345 6923 4379
rect 6647 4317 6681 4333
rect 6647 4133 6681 4149
rect 6957 4317 6991 4333
rect 6957 4133 6991 4149
rect 6715 4087 6731 4121
rect 6907 4087 6923 4121
rect 6647 4059 6681 4075
rect 6647 3875 6681 3891
rect 6957 4059 6991 4075
rect 6957 3875 6991 3891
rect 6715 3829 6731 3863
rect 6907 3829 6923 3863
rect 6647 3801 6681 3817
rect 6647 3617 6681 3633
rect 6957 3801 6991 3817
rect 6957 3617 6991 3633
rect 6715 3571 6731 3605
rect 6907 3571 6923 3605
rect 6647 3543 6681 3559
rect 6647 3359 6681 3375
rect 6957 3543 6991 3559
rect 6957 3359 6991 3375
rect 6715 3313 6731 3347
rect 6907 3313 6923 3347
rect 6647 3285 6681 3301
rect 6647 3101 6681 3117
rect 6957 3285 6991 3301
rect 6957 3101 6991 3117
rect 6715 3055 6731 3089
rect 6907 3055 6923 3089
rect 7094 2964 7141 8340
rect 6562 2963 7141 2964
rect 6343 2948 6473 2963
rect 6507 2948 7141 2963
rect 7175 2948 7233 8356
rect 7303 8068 8160 8070
rect 7301 8047 8160 8068
rect 7301 8013 7419 8047
rect 7793 8013 8160 8047
rect 7301 7992 8160 8013
rect 7301 7951 7369 7992
rect 7301 7423 7323 7951
rect 7357 7423 7369 7951
rect 7835 7951 8160 7992
rect 7502 7899 7518 7933
rect 7694 7899 7710 7933
rect 7425 7871 7459 7887
rect 7425 7487 7459 7503
rect 7753 7871 7787 7887
rect 7753 7487 7787 7503
rect 7502 7441 7518 7475
rect 7694 7441 7710 7475
rect 7301 7380 7369 7423
rect 7835 7423 7855 7951
rect 7889 7940 8160 7951
rect 7889 7423 7965 7940
rect 7835 7380 7965 7423
rect 7301 7361 7965 7380
rect 7301 7327 7419 7361
rect 7793 7327 7965 7361
rect 7301 7302 7965 7327
rect 7301 7301 7369 7302
rect 7307 6787 7383 6791
rect 7485 6787 7965 7302
rect 7307 6757 7965 6787
rect 7307 6723 7419 6757
rect 7793 6723 7965 6757
rect 7307 6702 7965 6723
rect 7307 6661 7383 6702
rect 7307 6133 7323 6661
rect 7357 6133 7383 6661
rect 7835 6661 7965 6702
rect 7502 6609 7518 6643
rect 7694 6609 7710 6643
rect 7425 6581 7459 6597
rect 7425 6197 7459 6213
rect 7753 6581 7787 6597
rect 7753 6197 7787 6213
rect 7502 6151 7518 6185
rect 7694 6151 7710 6185
rect 7307 6081 7383 6133
rect 7835 6133 7855 6661
rect 7889 6133 7965 6661
rect 7835 6081 7965 6133
rect 7307 6071 7965 6081
rect 7307 6037 7419 6071
rect 7793 6037 7965 6071
rect 7307 6001 7965 6037
rect 7473 5495 7965 6001
rect 7298 5467 7965 5495
rect 7298 5433 7419 5467
rect 7793 5433 7965 5467
rect 7298 5404 7965 5433
rect 7298 5371 7381 5404
rect 7298 4843 7323 5371
rect 7357 4843 7381 5371
rect 7834 5371 7965 5404
rect 7502 5319 7518 5353
rect 7694 5319 7710 5353
rect 7834 5308 7855 5371
rect 7425 5291 7459 5307
rect 7425 4907 7459 4923
rect 7753 5291 7787 5307
rect 7753 4907 7787 4923
rect 7502 4861 7518 4895
rect 7694 4861 7710 4895
rect 7298 4807 7381 4843
rect 7835 4843 7855 5308
rect 7889 4843 7965 5371
rect 7835 4808 7965 4843
rect 7834 4807 7965 4808
rect 7298 4781 7965 4807
rect 7298 4747 7419 4781
rect 7793 4747 7965 4781
rect 7298 4711 7965 4747
rect 7473 4203 7965 4711
rect 7309 4201 7965 4203
rect 6343 2922 7233 2948
rect 6343 2888 6533 2922
rect 7115 2888 7233 2922
rect 6343 2841 7233 2888
rect 7307 4164 7965 4201
rect 7307 4130 7407 4164
rect 7831 4130 7965 4164
rect 7307 4118 7965 4130
rect 7307 4104 7386 4118
rect 7307 2940 7347 4104
rect 7381 2940 7386 4104
rect 7835 4104 7965 4118
rect 7502 4029 7518 4063
rect 7694 4029 7710 4063
rect 7425 4001 7459 4017
rect 7425 3617 7459 3633
rect 7753 4001 7787 4017
rect 7753 3617 7787 3633
rect 7502 3571 7518 3605
rect 7694 3571 7710 3605
rect 7502 3448 7518 3482
rect 7694 3448 7710 3482
rect 7425 3420 7459 3436
rect 7425 3036 7459 3052
rect 7753 3420 7787 3436
rect 7753 3036 7787 3052
rect 7502 2990 7518 3024
rect 7694 2990 7710 3024
rect 7307 2935 7386 2940
rect 7835 2940 7857 4104
rect 7891 2945 7965 4104
rect 8104 4274 8160 7940
rect 17727 7384 19149 8938
rect 17726 7383 19149 7384
rect 17726 7349 17968 7383
rect 18724 7349 19149 7383
rect 17726 7347 19149 7349
rect 17726 7287 17937 7347
rect 17726 6159 17872 7287
rect 17906 6159 17937 7287
rect 18778 7287 19149 7347
rect 18042 7235 18058 7269
rect 18634 7235 18650 7269
rect 17974 7207 18008 7223
rect 17974 6223 18008 6239
rect 18684 7207 18718 7223
rect 18684 6223 18718 6239
rect 17726 6101 17937 6159
rect 18042 6177 18058 6211
rect 18634 6177 18650 6211
rect 18042 6101 18650 6177
rect 18778 6159 18786 7287
rect 18820 6159 19149 7287
rect 18778 6101 19149 6159
rect 17726 6097 19149 6101
rect 17726 6063 17968 6097
rect 18724 6063 19149 6097
rect 17726 5871 19149 6063
rect 17724 5667 19149 5871
rect 17724 5573 17832 5667
rect 18385 5596 19149 5667
rect 19183 8925 24536 8938
rect 19183 5596 19203 8925
rect 19431 8832 19447 8866
rect 21815 8832 21831 8866
rect 21889 8832 21905 8866
rect 24273 8832 24289 8866
rect 19385 8782 19419 8798
rect 19385 7590 19419 7606
rect 21843 8782 21877 8798
rect 21843 7590 21877 7606
rect 24301 8782 24335 8798
rect 24301 7590 24335 7606
rect 19431 7522 19447 7556
rect 21815 7522 21831 7556
rect 21889 7522 21905 7556
rect 24273 7522 24289 7556
rect 19430 6957 19446 6991
rect 21814 6957 21830 6991
rect 21888 6957 21904 6991
rect 24272 6957 24288 6991
rect 19384 6907 19418 6923
rect 19384 5715 19418 5731
rect 21842 6907 21876 6923
rect 21842 5715 21876 5731
rect 24300 6907 24334 6923
rect 24300 5715 24334 5731
rect 19430 5647 19446 5681
rect 21814 5647 21830 5681
rect 21888 5647 21904 5681
rect 24272 5647 24288 5681
rect 18385 5591 19203 5596
rect 24526 5596 24536 8925
rect 24570 5596 24876 8938
rect 24526 5591 24876 5596
rect 18385 5573 24876 5591
rect 17724 5570 24876 5573
rect 17724 5536 19209 5570
rect 24510 5536 24876 5570
rect 17724 5432 24876 5536
rect 17724 5343 17834 5432
rect 24768 5343 24876 5432
rect 17724 5281 24876 5343
rect 8104 2945 8161 4274
rect 7891 2940 8161 2945
rect 7835 2935 8161 2940
rect 7307 2914 8161 2935
rect 7307 2880 7407 2914
rect 7831 2880 8161 2914
rect 7307 2832 8161 2880
rect 7307 2831 7851 2832
<< viali >>
rect 3401 30801 11199 30890
rect 3728 30499 7296 30533
rect 7386 30499 10954 30533
rect 3666 30104 3700 30440
rect 7324 30104 7358 30440
rect 10982 30104 11016 30440
rect 3728 30011 7296 30045
rect 7386 30011 10954 30045
rect 3666 29616 3700 29952
rect 7324 29616 7358 29952
rect 10982 29616 11016 29952
rect 3728 29523 7296 29557
rect 7386 29523 10954 29557
rect 11800 32942 14392 33012
rect 11800 32908 11934 32942
rect 11934 32908 14214 32942
rect 14214 32908 14392 32942
rect 11800 32882 14392 32908
rect 11800 29401 11874 32882
rect 11874 29401 11908 32882
rect 11908 32809 14240 32882
rect 14240 32809 14274 32882
rect 14274 32809 14392 32882
rect 11908 29401 11965 32809
rect 12200 32575 12548 32609
rect 12638 32575 12986 32609
rect 13076 32575 13424 32609
rect 13514 32575 13862 32609
rect 12138 29540 12172 32516
rect 12576 29540 12610 32516
rect 13014 29540 13048 32516
rect 13452 29540 13486 32516
rect 13890 29540 13924 32516
rect 14180 29750 14240 32230
rect 14240 29750 14274 32230
rect 14274 29750 14322 32230
rect 12200 29447 12548 29481
rect 12638 29447 12986 29481
rect 13076 29447 13424 29481
rect 13514 29447 13862 29481
rect 3549 27021 4125 27055
rect 3465 26025 3499 26993
rect 4175 26025 4209 26993
rect 3549 25963 4125 25997
rect 3323 25359 3876 25453
rect 4938 28618 7306 28652
rect 7396 28618 9764 28652
rect 4876 27392 4910 28568
rect 7334 27392 7368 28568
rect 9792 27392 9826 28568
rect 4938 27308 7306 27342
rect 7396 27308 9764 27342
rect 4937 26743 7305 26777
rect 7395 26743 9763 26777
rect 4875 25517 4909 26693
rect 7333 25517 7367 26693
rect 9791 25517 9825 26693
rect 4937 25433 7305 25467
rect 7395 25433 9763 25467
rect 12200 28598 12548 28632
rect 12638 28598 12986 28632
rect 13076 28598 13424 28632
rect 13514 28598 13862 28632
rect 11817 25407 11874 28583
rect 11816 25347 11874 25407
rect 11874 25347 11908 28583
rect 11908 25374 11965 28583
rect 12138 25563 12172 28539
rect 12576 25563 12610 28539
rect 13014 25563 13048 28539
rect 13452 25563 13486 28539
rect 13890 25563 13924 28539
rect 14196 25517 14240 27997
rect 14240 25517 14274 27997
rect 14274 27499 14338 27997
rect 25403 28157 25662 28158
rect 20700 27858 25662 28157
rect 20700 27824 20855 27858
rect 20855 27824 25541 27858
rect 25541 27824 25662 27858
rect 20700 27798 25662 27824
rect 20700 27792 20795 27798
rect 14274 27498 19128 27499
rect 14274 27207 19138 27498
rect 14274 25517 14338 27207
rect 12200 25470 12548 25504
rect 12638 25470 12986 25504
rect 13076 25470 13424 25504
rect 13514 25470 13862 25504
rect 11908 25347 14240 25374
rect 14240 25347 14274 25374
rect 14274 25347 14381 25374
rect 11816 25321 14381 25347
rect 11816 25287 11934 25321
rect 11934 25287 14214 25321
rect 14214 25287 14381 25321
rect 11816 25231 14381 25287
rect 11929 25230 14381 25231
rect 3325 25129 10259 25218
rect 16600 25451 16833 27207
rect 17029 27044 17357 27078
rect 17447 27044 17775 27078
rect 17865 27044 18193 27078
rect 18283 27044 18611 27078
rect 16967 25609 17001 26985
rect 17385 25609 17419 26985
rect 17803 25609 17837 26985
rect 18221 25609 18255 26985
rect 18639 25609 18673 26985
rect 17029 25516 17357 25550
rect 17447 25516 17775 25550
rect 17865 25516 18193 25550
rect 18283 25516 18611 25550
rect 18851 25691 19138 27207
rect 20762 25585 20795 27792
rect 20795 25585 20829 27798
rect 20829 27793 25567 27798
rect 20829 27792 25504 27793
rect 20829 25590 20879 27792
rect 21122 27589 22090 27623
rect 22180 27589 23148 27623
rect 23238 27589 24206 27623
rect 24296 27589 25264 27623
rect 21060 27054 21094 27530
rect 22118 27054 22152 27530
rect 23176 27054 23210 27530
rect 24234 27054 24268 27530
rect 25292 27054 25326 27530
rect 21122 26961 22090 26995
rect 22180 26961 23148 26995
rect 23238 26961 24206 26995
rect 24296 26961 25264 26995
rect 25546 26979 25567 27793
rect 25567 26979 25601 27798
rect 25601 27793 25662 27798
rect 25601 26979 25643 27793
rect 21122 26427 22090 26461
rect 22180 26427 23148 26461
rect 23238 26427 24206 26461
rect 24296 26427 25264 26461
rect 21060 25892 21094 26368
rect 22118 25892 22152 26368
rect 23176 25892 23210 26368
rect 24234 25892 24268 26368
rect 25292 25892 25326 26368
rect 21122 25799 22090 25833
rect 22180 25799 23148 25833
rect 23238 25799 24206 25833
rect 24296 25799 25264 25833
rect 20829 25585 25311 25590
rect 20762 25559 25311 25585
rect 20762 25525 20855 25559
rect 20855 25525 25311 25559
rect 20762 25500 25311 25525
rect 20797 25493 25311 25500
rect 16600 25448 18748 25451
rect 16600 25414 16949 25448
rect 16949 25414 18691 25448
rect 18691 25414 18748 25448
rect 16600 25217 18748 25414
rect 16685 25215 18748 25217
rect 22120 25311 24269 25360
rect 22120 25277 22195 25311
rect 22195 25277 24177 25311
rect 24177 25277 24269 25311
rect 22120 25257 24269 25277
rect 22120 25251 22178 25257
rect 11872 24889 12019 24892
rect 19698 24889 19814 24929
rect 11872 24855 11986 24889
rect 11986 24884 12019 24889
rect 11986 24883 12148 24884
rect 19698 24883 19814 24889
rect 11986 24855 19814 24883
rect 11872 24829 19814 24855
rect 11872 23606 11926 24829
rect 11926 23606 11960 24829
rect 11960 24780 19814 24829
rect 11960 23606 12019 24780
rect 19698 24768 19814 24780
rect 12210 24563 14058 24597
rect 14148 24563 15996 24597
rect 16086 24563 17934 24597
rect 18024 24563 19872 24597
rect 12148 24237 12182 24513
rect 14086 24237 14120 24513
rect 16024 24237 16058 24513
rect 17962 24237 17996 24513
rect 19900 24237 19934 24513
rect 12210 24153 14058 24187
rect 14148 24153 15996 24187
rect 16086 24153 17934 24187
rect 18024 24153 19872 24187
rect 12148 23827 12182 24103
rect 14086 23827 14120 24103
rect 16024 23827 16058 24103
rect 17962 23827 17996 24103
rect 19900 23827 19934 24103
rect 12210 23743 14058 23777
rect 14148 23743 15996 23777
rect 16086 23743 17934 23777
rect 18024 23743 19872 23777
rect 11872 23590 12019 23606
rect 11872 23589 12113 23590
rect 11872 23580 19791 23589
rect 11872 23546 11986 23580
rect 11986 23546 19791 23580
rect 11872 23392 19791 23546
rect 22120 24719 22135 25251
rect 22135 24719 22169 25251
rect 22169 24719 22178 25251
rect 24193 25251 24269 25257
rect 22307 25133 22675 25167
rect 22765 25133 23133 25167
rect 23223 25133 23591 25167
rect 23681 25133 24049 25167
rect 22245 24507 22279 25083
rect 22703 24507 22737 25083
rect 23161 24507 23195 25083
rect 23619 24507 23653 25083
rect 24077 24507 24111 25083
rect 22307 24423 22675 24457
rect 22765 24423 23133 24457
rect 23223 24423 23591 24457
rect 23681 24423 24049 24457
rect 22307 23926 22675 23960
rect 22765 23926 23133 23960
rect 23223 23926 23591 23960
rect 23681 23926 24049 23960
rect 22111 23133 22135 23683
rect 22135 23133 22169 23683
rect 22169 23133 22185 23683
rect 22245 23300 22279 23876
rect 22703 23300 22737 23876
rect 23161 23300 23195 23876
rect 23619 23300 23653 23876
rect 24077 23300 24111 23876
rect 22307 23216 22675 23250
rect 22765 23216 23133 23250
rect 23223 23216 23591 23250
rect 23681 23216 24049 23250
rect 22111 23052 22185 23133
rect 24193 23133 24203 25251
rect 24203 23133 24237 25251
rect 24237 23133 24269 25251
rect 25207 25064 25311 25493
rect 25207 24370 25279 25064
rect 25279 24370 25311 25064
rect 25455 25024 25493 25058
rect 25393 24469 25427 24965
rect 25521 24469 25555 24965
rect 25455 24376 25493 24410
rect 25207 24334 25311 24370
rect 25811 25024 25849 25058
rect 25749 24469 25783 24965
rect 25877 24469 25911 24965
rect 25811 24376 25849 24410
rect 25477 24010 25511 24044
rect 25833 24010 25867 24044
rect 25433 23784 25467 23960
rect 25521 23784 25555 23960
rect 25789 23784 25823 23960
rect 25877 23784 25911 23960
rect 25477 23700 25511 23734
rect 25833 23700 25867 23734
rect 24611 23228 25989 23500
rect 24193 23052 24269 23133
rect 24611 23052 24731 23228
rect 22066 22882 24731 23052
rect 24907 22962 25304 23000
rect 25546 22962 25943 23000
rect 12053 21654 12227 21700
rect 14994 21654 15106 21656
rect 12053 15198 12190 21654
rect 12190 15198 12224 21654
rect 12224 15198 12227 21654
rect 12478 21536 13254 21570
rect 13959 21536 14735 21570
rect 12394 21340 12428 21508
rect 13304 21340 13338 21508
rect 13875 21340 13909 21508
rect 14785 21340 14819 21508
rect 12478 21278 13254 21312
rect 13959 21278 14735 21312
rect 12394 21082 12428 21250
rect 13304 21082 13338 21250
rect 13875 21082 13909 21250
rect 14785 21082 14819 21250
rect 12478 21020 13254 21054
rect 13959 21020 14735 21054
rect 12394 20824 12428 20992
rect 13304 20824 13338 20992
rect 13875 20824 13909 20992
rect 14785 20824 14819 20992
rect 12478 20762 13254 20796
rect 13959 20762 14735 20796
rect 12394 20566 12428 20734
rect 13304 20566 13338 20734
rect 13875 20566 13909 20734
rect 14785 20566 14819 20734
rect 12478 20504 13254 20538
rect 13959 20504 14735 20538
rect 12394 20308 12428 20476
rect 13304 20308 13338 20476
rect 13875 20308 13909 20476
rect 14785 20308 14819 20476
rect 12478 20246 13254 20280
rect 13959 20246 14735 20280
rect 12394 20050 12428 20218
rect 13304 20050 13338 20218
rect 13875 20050 13909 20218
rect 14785 20050 14819 20218
rect 12478 19988 13254 20022
rect 13959 19988 14735 20022
rect 12394 19792 12428 19960
rect 13304 19792 13338 19960
rect 13875 19792 13909 19960
rect 14785 19792 14819 19960
rect 12478 19730 13254 19764
rect 13959 19730 14735 19764
rect 12394 19534 12428 19702
rect 13304 19534 13338 19702
rect 13875 19534 13909 19702
rect 14785 19534 14819 19702
rect 12478 19472 13254 19506
rect 13959 19472 14735 19506
rect 12394 19276 12428 19444
rect 13304 19276 13338 19444
rect 13875 19276 13909 19444
rect 14785 19276 14819 19444
rect 12478 19214 13254 19248
rect 13959 19214 14735 19248
rect 12394 19018 12428 19186
rect 13304 19018 13338 19186
rect 13875 19018 13909 19186
rect 14785 19018 14819 19186
rect 12478 18956 13254 18990
rect 13959 18956 14735 18990
rect 12394 18760 12428 18928
rect 13304 18760 13338 18928
rect 13875 18760 13909 18928
rect 14785 18760 14819 18928
rect 12478 18698 13254 18732
rect 13959 18698 14735 18732
rect 12394 18502 12428 18670
rect 13304 18502 13338 18670
rect 13875 18502 13909 18670
rect 14785 18502 14819 18670
rect 12478 18440 13254 18474
rect 13959 18440 14735 18474
rect 12394 18244 12428 18412
rect 13304 18244 13338 18412
rect 13875 18244 13909 18412
rect 14785 18244 14819 18412
rect 12478 18182 13254 18216
rect 13959 18182 14735 18216
rect 12394 17986 12428 18154
rect 13304 17986 13338 18154
rect 13875 17986 13909 18154
rect 14785 17986 14819 18154
rect 12478 17924 13254 17958
rect 13959 17924 14735 17958
rect 12394 17728 12428 17896
rect 13304 17728 13338 17896
rect 13875 17728 13909 17896
rect 14785 17728 14819 17896
rect 12478 17666 13254 17700
rect 13959 17666 14735 17700
rect 12394 17470 12428 17638
rect 13304 17470 13338 17638
rect 13875 17470 13909 17638
rect 14785 17470 14819 17638
rect 12478 17408 13254 17442
rect 13959 17408 14735 17442
rect 12394 17212 12428 17380
rect 13304 17212 13338 17380
rect 13875 17212 13909 17380
rect 14785 17212 14819 17380
rect 12478 17150 13254 17184
rect 13959 17150 14735 17184
rect 12394 16954 12428 17122
rect 13304 16954 13338 17122
rect 13875 16954 13909 17122
rect 14785 16954 14819 17122
rect 12478 16892 13254 16926
rect 13959 16892 14735 16926
rect 12394 16696 12428 16864
rect 13304 16696 13338 16864
rect 13875 16696 13909 16864
rect 14785 16696 14819 16864
rect 12478 16634 13254 16668
rect 13959 16634 14735 16668
rect 12394 16438 12428 16606
rect 13304 16438 13338 16606
rect 13875 16438 13909 16606
rect 14785 16438 14819 16606
rect 12478 16376 13254 16410
rect 13959 16376 14735 16410
rect 12394 16180 12428 16348
rect 13304 16180 13338 16348
rect 13875 16180 13909 16348
rect 14785 16180 14819 16348
rect 12478 16118 13254 16152
rect 13959 16118 14735 16152
rect 12394 15922 12428 16090
rect 13304 15922 13338 16090
rect 13875 15922 13909 16090
rect 14785 15922 14819 16090
rect 12478 15860 13254 15894
rect 13959 15860 14735 15894
rect 12394 15664 12428 15832
rect 13304 15664 13338 15832
rect 13875 15664 13909 15832
rect 14785 15664 14819 15832
rect 12478 15602 13254 15636
rect 13959 15602 14735 15636
rect 12394 15406 12428 15574
rect 13304 15406 13338 15574
rect 13875 15406 13909 15574
rect 14785 15406 14819 15574
rect 12478 15344 13254 15378
rect 13959 15344 14735 15378
rect 14994 15315 15019 21654
rect 15019 15315 15106 21654
rect 15736 17074 15838 22467
rect 15838 17074 15872 22467
rect 15872 17074 15927 22467
rect 16096 22341 16272 22375
rect 16012 22145 16046 22313
rect 16322 22145 16356 22313
rect 16096 22083 16272 22117
rect 16012 21887 16046 22055
rect 16322 21887 16356 22055
rect 16096 21825 16272 21859
rect 16012 21629 16046 21797
rect 16322 21629 16356 21797
rect 16096 21567 16272 21601
rect 16012 21371 16046 21539
rect 16322 21371 16356 21539
rect 16096 21309 16272 21343
rect 16012 21113 16046 21281
rect 16322 21113 16356 21281
rect 16096 21051 16272 21085
rect 16012 20855 16046 21023
rect 16322 20855 16356 21023
rect 16096 20793 16272 20827
rect 16012 20597 16046 20765
rect 16322 20597 16356 20765
rect 16096 20535 16272 20569
rect 16012 20339 16046 20507
rect 16322 20339 16356 20507
rect 16096 20277 16272 20311
rect 16012 20081 16046 20249
rect 16322 20081 16356 20249
rect 16096 20019 16272 20053
rect 16012 19823 16046 19991
rect 16322 19823 16356 19991
rect 16096 19761 16272 19795
rect 16012 19565 16046 19733
rect 16322 19565 16356 19733
rect 16096 19503 16272 19537
rect 16012 19307 16046 19475
rect 16322 19307 16356 19475
rect 16096 19245 16272 19279
rect 16012 19049 16046 19217
rect 16322 19049 16356 19217
rect 16096 18987 16272 19021
rect 16012 18791 16046 18959
rect 16322 18791 16356 18959
rect 16096 18729 16272 18763
rect 16012 18533 16046 18701
rect 16322 18533 16356 18701
rect 16096 18471 16272 18505
rect 16012 18275 16046 18443
rect 16322 18275 16356 18443
rect 16096 18213 16272 18247
rect 16012 18017 16046 18185
rect 16322 18017 16356 18185
rect 16096 17955 16272 17989
rect 16012 17759 16046 17927
rect 16322 17759 16356 17927
rect 16096 17697 16272 17731
rect 16012 17501 16046 17669
rect 16322 17501 16356 17669
rect 16096 17439 16272 17473
rect 16012 17243 16046 17411
rect 16322 17243 16356 17411
rect 16096 17181 16272 17215
rect 16883 22406 17059 22440
rect 16790 22010 16824 22378
rect 17118 22010 17152 22378
rect 16883 21948 17059 21982
rect 16883 21825 17059 21859
rect 16790 21429 16824 21797
rect 17118 21429 17152 21797
rect 16883 21367 17059 21401
rect 16883 20535 17059 20569
rect 16790 20139 16824 20507
rect 17118 20139 17152 20507
rect 16883 20077 17059 20111
rect 16883 19245 17059 19279
rect 16790 18849 16824 19217
rect 17118 18849 17152 19217
rect 16883 18787 17059 18821
rect 16883 17955 17059 17989
rect 16790 17559 16824 17927
rect 17118 17559 17152 17927
rect 16883 17497 17059 17531
rect 17330 17490 17469 22485
rect 22066 21866 22404 22882
rect 22666 22716 23742 22750
rect 22582 22420 22616 22688
rect 23792 22420 23826 22688
rect 22666 22358 23742 22392
rect 22582 22062 22616 22330
rect 23792 22062 23826 22330
rect 22666 22000 23742 22034
rect 23955 21866 24166 22882
rect 22066 21627 24166 21866
rect 22066 21625 22293 21627
rect 23955 21616 24166 21627
rect 15736 17060 15927 17074
rect 17251 16941 17351 17028
rect 16883 16867 17059 16901
rect 17216 16899 17351 16941
rect 16790 16671 16824 16839
rect 17118 16671 17152 16839
rect 15334 16210 16377 16316
rect 15334 16208 15494 16210
rect 15494 16208 15528 16210
rect 15528 16208 15584 16210
rect 15584 16208 15618 16210
rect 15618 16208 15674 16210
rect 15674 16208 15708 16210
rect 15708 16208 15764 16210
rect 15764 16208 15798 16210
rect 15798 16208 15854 16210
rect 15854 16208 15888 16210
rect 15888 16208 15944 16210
rect 15944 16208 15978 16210
rect 15978 16208 16034 16210
rect 16034 16208 16068 16210
rect 16068 16208 16124 16210
rect 16124 16208 16158 16210
rect 16158 16208 16214 16210
rect 16214 16208 16248 16210
rect 16248 16208 16377 16210
rect 15155 15307 15251 15834
rect 15620 16002 15626 16008
rect 15626 16002 15654 16008
rect 15620 15974 15654 16002
rect 15720 15974 15754 16008
rect 15820 15974 15854 16008
rect 15920 16002 15952 16008
rect 15952 16002 15954 16008
rect 16020 16002 16042 16008
rect 16042 16002 16054 16008
rect 16120 16002 16132 16008
rect 16132 16002 16154 16008
rect 15920 15974 15954 16002
rect 16020 15974 16054 16002
rect 16120 15974 16154 16002
rect 15620 15874 15654 15908
rect 15720 15874 15754 15908
rect 15820 15874 15854 15908
rect 15920 15874 15954 15908
rect 16020 15874 16054 15908
rect 16120 15874 16154 15908
rect 15620 15774 15654 15808
rect 15720 15774 15754 15808
rect 15820 15774 15854 15808
rect 15920 15774 15954 15808
rect 16020 15774 16054 15808
rect 16120 15774 16154 15808
rect 15620 15676 15654 15708
rect 15620 15674 15626 15676
rect 15626 15674 15654 15676
rect 15720 15674 15754 15708
rect 15820 15674 15854 15708
rect 15920 15676 15954 15708
rect 16020 15676 16054 15708
rect 16120 15676 16154 15708
rect 15920 15674 15952 15676
rect 15952 15674 15954 15676
rect 16020 15674 16042 15676
rect 16042 15674 16054 15676
rect 16120 15674 16132 15676
rect 16132 15674 16154 15676
rect 15620 15586 15654 15608
rect 15620 15574 15626 15586
rect 15626 15574 15654 15586
rect 15720 15574 15754 15608
rect 15820 15574 15854 15608
rect 15920 15586 15954 15608
rect 16020 15586 16054 15608
rect 16120 15586 16154 15608
rect 15920 15574 15952 15586
rect 15952 15574 15954 15586
rect 16020 15574 16042 15586
rect 16042 15574 16054 15586
rect 16120 15574 16132 15586
rect 16132 15574 16154 15586
rect 15620 15496 15654 15508
rect 15620 15474 15626 15496
rect 15626 15474 15654 15496
rect 15720 15474 15754 15508
rect 15820 15474 15854 15508
rect 15920 15496 15954 15508
rect 16020 15496 16054 15508
rect 16120 15496 16154 15508
rect 15920 15474 15952 15496
rect 15952 15474 15954 15496
rect 16020 15474 16042 15496
rect 16042 15474 16054 15496
rect 16120 15474 16132 15496
rect 16132 15474 16154 15496
rect 16344 16078 16492 16083
rect 16344 16044 16458 16078
rect 16458 16044 16492 16078
rect 16344 15988 16492 16044
rect 16344 15954 16458 15988
rect 16458 15954 16492 15988
rect 16344 15898 16492 15954
rect 16344 15864 16458 15898
rect 16458 15864 16492 15898
rect 16344 15808 16492 15864
rect 16344 15774 16458 15808
rect 16458 15774 16492 15808
rect 16344 15718 16492 15774
rect 16344 15684 16458 15718
rect 16458 15684 16492 15718
rect 16344 15628 16492 15684
rect 16344 15594 16458 15628
rect 16458 15594 16492 15628
rect 16344 15538 16492 15594
rect 16344 15504 16458 15538
rect 16458 15504 16492 15538
rect 16344 15448 16492 15504
rect 16344 15414 16458 15448
rect 16458 15414 16492 15448
rect 16344 15358 16492 15414
rect 16344 15324 16458 15358
rect 16458 15324 16492 15358
rect 12053 15122 12227 15198
rect 12309 15172 12461 15179
rect 13299 15172 13447 15179
rect 15767 15172 16246 15281
rect 16344 15268 16492 15324
rect 16344 15258 16458 15268
rect 16458 15258 16492 15268
rect 12309 15138 12461 15172
rect 13299 15138 13447 15172
rect 15767 15161 15778 15172
rect 15778 15161 15834 15172
rect 15834 15161 15868 15172
rect 15868 15161 15924 15172
rect 15924 15161 15958 15172
rect 15958 15161 16014 15172
rect 16014 15161 16048 15172
rect 16048 15161 16104 15172
rect 16104 15161 16138 15172
rect 16138 15161 16194 15172
rect 16194 15161 16228 15172
rect 16228 15161 16246 15172
rect 12309 15125 12461 15138
rect 13299 15125 13447 15138
rect 16883 16609 17059 16643
rect 16790 16413 16824 16581
rect 17118 16413 17152 16581
rect 16883 16351 17059 16385
rect 16883 16142 16959 16176
rect 16790 15746 16824 16114
rect 17018 15746 17052 16114
rect 16883 15684 16959 15718
rect 16790 15288 16824 15656
rect 17018 15288 17052 15656
rect 17216 16042 17247 16899
rect 17247 16042 17351 16899
rect 16883 15226 16959 15260
rect 17218 15224 17247 16042
rect 17247 15224 17350 16042
rect 17218 15049 17350 15224
rect 17429 15050 17577 17029
rect 17910 11015 25708 11104
rect 2688 10331 2862 10407
rect 2944 10391 3096 10404
rect 3934 10391 4082 10404
rect 2944 10357 3096 10391
rect 3934 10357 4082 10391
rect 6402 10357 6413 10368
rect 6413 10357 6469 10368
rect 6469 10357 6503 10368
rect 6503 10357 6559 10368
rect 6559 10357 6593 10368
rect 6593 10357 6649 10368
rect 6649 10357 6683 10368
rect 6683 10357 6739 10368
rect 6739 10357 6773 10368
rect 6773 10357 6829 10368
rect 6829 10357 6863 10368
rect 6863 10357 6881 10368
rect 2944 10350 3096 10357
rect 3934 10350 4082 10357
rect 2688 3875 2825 10331
rect 2825 3875 2859 10331
rect 2859 3875 2862 10331
rect 3113 10151 3889 10185
rect 4594 10151 5370 10185
rect 6402 10248 6881 10357
rect 6979 10261 7093 10271
rect 7093 10261 7127 10271
rect 3029 9955 3063 10123
rect 3939 9955 3973 10123
rect 4510 9955 4544 10123
rect 5420 9955 5454 10123
rect 3113 9893 3889 9927
rect 4594 9893 5370 9927
rect 3029 9697 3063 9865
rect 3939 9697 3973 9865
rect 4510 9697 4544 9865
rect 5420 9697 5454 9865
rect 3113 9635 3889 9669
rect 4594 9635 5370 9669
rect 3029 9439 3063 9607
rect 3939 9439 3973 9607
rect 4510 9439 4544 9607
rect 5420 9439 5454 9607
rect 3113 9377 3889 9411
rect 4594 9377 5370 9411
rect 3029 9181 3063 9349
rect 3939 9181 3973 9349
rect 4510 9181 4544 9349
rect 5420 9181 5454 9349
rect 3113 9119 3889 9153
rect 4594 9119 5370 9153
rect 3029 8923 3063 9091
rect 3939 8923 3973 9091
rect 4510 8923 4544 9091
rect 5420 8923 5454 9091
rect 3113 8861 3889 8895
rect 4594 8861 5370 8895
rect 3029 8665 3063 8833
rect 3939 8665 3973 8833
rect 4510 8665 4544 8833
rect 5420 8665 5454 8833
rect 3113 8603 3889 8637
rect 4594 8603 5370 8637
rect 3029 8407 3063 8575
rect 3939 8407 3973 8575
rect 4510 8407 4544 8575
rect 5420 8407 5454 8575
rect 3113 8345 3889 8379
rect 4594 8345 5370 8379
rect 3029 8149 3063 8317
rect 3939 8149 3973 8317
rect 4510 8149 4544 8317
rect 5420 8149 5454 8317
rect 3113 8087 3889 8121
rect 4594 8087 5370 8121
rect 3029 7891 3063 8059
rect 3939 7891 3973 8059
rect 4510 7891 4544 8059
rect 5420 7891 5454 8059
rect 3113 7829 3889 7863
rect 4594 7829 5370 7863
rect 3029 7633 3063 7801
rect 3939 7633 3973 7801
rect 4510 7633 4544 7801
rect 5420 7633 5454 7801
rect 3113 7571 3889 7605
rect 4594 7571 5370 7605
rect 3029 7375 3063 7543
rect 3939 7375 3973 7543
rect 4510 7375 4544 7543
rect 5420 7375 5454 7543
rect 3113 7313 3889 7347
rect 4594 7313 5370 7347
rect 3029 7117 3063 7285
rect 3939 7117 3973 7285
rect 4510 7117 4544 7285
rect 5420 7117 5454 7285
rect 3113 7055 3889 7089
rect 4594 7055 5370 7089
rect 3029 6859 3063 7027
rect 3939 6859 3973 7027
rect 4510 6859 4544 7027
rect 5420 6859 5454 7027
rect 3113 6797 3889 6831
rect 4594 6797 5370 6831
rect 3029 6601 3063 6769
rect 3939 6601 3973 6769
rect 4510 6601 4544 6769
rect 5420 6601 5454 6769
rect 3113 6539 3889 6573
rect 4594 6539 5370 6573
rect 3029 6343 3063 6511
rect 3939 6343 3973 6511
rect 4510 6343 4544 6511
rect 5420 6343 5454 6511
rect 3113 6281 3889 6315
rect 4594 6281 5370 6315
rect 3029 6085 3063 6253
rect 3939 6085 3973 6253
rect 4510 6085 4544 6253
rect 5420 6085 5454 6253
rect 3113 6023 3889 6057
rect 4594 6023 5370 6057
rect 3029 5827 3063 5995
rect 3939 5827 3973 5995
rect 4510 5827 4544 5995
rect 5420 5827 5454 5995
rect 3113 5765 3889 5799
rect 4594 5765 5370 5799
rect 3029 5569 3063 5737
rect 3939 5569 3973 5737
rect 4510 5569 4544 5737
rect 5420 5569 5454 5737
rect 3113 5507 3889 5541
rect 4594 5507 5370 5541
rect 3029 5311 3063 5479
rect 3939 5311 3973 5479
rect 4510 5311 4544 5479
rect 5420 5311 5454 5479
rect 3113 5249 3889 5283
rect 4594 5249 5370 5283
rect 3029 5053 3063 5221
rect 3939 5053 3973 5221
rect 4510 5053 4544 5221
rect 5420 5053 5454 5221
rect 3113 4991 3889 5025
rect 4594 4991 5370 5025
rect 3029 4795 3063 4963
rect 3939 4795 3973 4963
rect 4510 4795 4544 4963
rect 5420 4795 5454 4963
rect 3113 4733 3889 4767
rect 4594 4733 5370 4767
rect 3029 4537 3063 4705
rect 3939 4537 3973 4705
rect 4510 4537 4544 4705
rect 5420 4537 5454 4705
rect 3113 4475 3889 4509
rect 4594 4475 5370 4509
rect 3029 4279 3063 4447
rect 3939 4279 3973 4447
rect 4510 4279 4544 4447
rect 5420 4279 5454 4447
rect 3113 4217 3889 4251
rect 4594 4217 5370 4251
rect 3029 4021 3063 4189
rect 3939 4021 3973 4189
rect 4510 4021 4544 4189
rect 5420 4021 5454 4189
rect 3113 3959 3889 3993
rect 4594 3959 5370 3993
rect 5629 3875 5654 10214
rect 5654 3875 5741 10214
rect 5790 9695 5886 10222
rect 6979 10205 7127 10261
rect 6979 10171 7093 10205
rect 7093 10171 7127 10205
rect 6255 10033 6261 10055
rect 6261 10033 6289 10055
rect 6255 10021 6289 10033
rect 6355 10021 6389 10055
rect 6455 10021 6489 10055
rect 6555 10033 6587 10055
rect 6587 10033 6589 10055
rect 6655 10033 6677 10055
rect 6677 10033 6689 10055
rect 6755 10033 6767 10055
rect 6767 10033 6789 10055
rect 6555 10021 6589 10033
rect 6655 10021 6689 10033
rect 6755 10021 6789 10033
rect 6255 9943 6261 9955
rect 6261 9943 6289 9955
rect 6255 9921 6289 9943
rect 6355 9921 6389 9955
rect 6455 9921 6489 9955
rect 6555 9943 6587 9955
rect 6587 9943 6589 9955
rect 6655 9943 6677 9955
rect 6677 9943 6689 9955
rect 6755 9943 6767 9955
rect 6767 9943 6789 9955
rect 6555 9921 6589 9943
rect 6655 9921 6689 9943
rect 6755 9921 6789 9943
rect 6255 9853 6261 9855
rect 6261 9853 6289 9855
rect 6255 9821 6289 9853
rect 6355 9821 6389 9855
rect 6455 9821 6489 9855
rect 6555 9853 6587 9855
rect 6587 9853 6589 9855
rect 6655 9853 6677 9855
rect 6677 9853 6689 9855
rect 6755 9853 6767 9855
rect 6767 9853 6789 9855
rect 6555 9821 6589 9853
rect 6655 9821 6689 9853
rect 6755 9821 6789 9853
rect 6255 9721 6289 9755
rect 6355 9721 6389 9755
rect 6455 9721 6489 9755
rect 6555 9721 6589 9755
rect 6655 9721 6689 9755
rect 6755 9721 6789 9755
rect 6255 9621 6289 9655
rect 6355 9621 6389 9655
rect 6455 9621 6489 9655
rect 6555 9621 6589 9655
rect 6655 9621 6689 9655
rect 6755 9621 6789 9655
rect 6255 9527 6289 9555
rect 6255 9521 6261 9527
rect 6261 9521 6289 9527
rect 6355 9521 6389 9555
rect 6455 9521 6489 9555
rect 6555 9527 6589 9555
rect 6655 9527 6689 9555
rect 6755 9527 6789 9555
rect 6555 9521 6587 9527
rect 6587 9521 6589 9527
rect 6655 9521 6677 9527
rect 6677 9521 6689 9527
rect 6755 9521 6767 9527
rect 6767 9521 6789 9527
rect 6979 10115 7127 10171
rect 6979 10081 7093 10115
rect 7093 10081 7127 10115
rect 6979 10025 7127 10081
rect 6979 9991 7093 10025
rect 7093 9991 7127 10025
rect 6979 9935 7127 9991
rect 6979 9901 7093 9935
rect 7093 9901 7127 9935
rect 6979 9845 7127 9901
rect 6979 9811 7093 9845
rect 7093 9811 7127 9845
rect 6979 9755 7127 9811
rect 6979 9721 7093 9755
rect 7093 9721 7127 9755
rect 6979 9665 7127 9721
rect 6979 9631 7093 9665
rect 7093 9631 7127 9665
rect 6979 9575 7127 9631
rect 6979 9541 7093 9575
rect 7093 9541 7127 9575
rect 6979 9485 7127 9541
rect 6979 9451 7093 9485
rect 7093 9451 7127 9485
rect 6979 9446 7127 9451
rect 5969 9319 6129 9321
rect 6129 9319 6163 9321
rect 6163 9319 6219 9321
rect 6219 9319 6253 9321
rect 6253 9319 6309 9321
rect 6309 9319 6343 9321
rect 6343 9319 6399 9321
rect 6399 9319 6433 9321
rect 6433 9319 6489 9321
rect 6489 9319 6523 9321
rect 6523 9319 6579 9321
rect 6579 9319 6613 9321
rect 6613 9319 6669 9321
rect 6669 9319 6703 9321
rect 6703 9319 6759 9321
rect 6759 9319 6793 9321
rect 6793 9319 6849 9321
rect 6849 9319 6883 9321
rect 6883 9319 7012 9321
rect 5969 9213 7012 9319
rect 7853 10305 7985 10480
rect 7518 10269 7594 10303
rect 7425 9873 7459 10241
rect 7653 9873 7687 10241
rect 7518 9811 7594 9845
rect 7425 9415 7459 9783
rect 7653 9415 7687 9783
rect 7518 9353 7594 9387
rect 7853 9487 7882 10305
rect 7882 9487 7985 10305
rect 7518 9144 7694 9178
rect 7425 8948 7459 9116
rect 7753 8948 7787 9116
rect 7518 8886 7694 8920
rect 7425 8690 7459 8858
rect 7753 8690 7787 8858
rect 7518 8628 7694 8662
rect 7851 8630 7882 9487
rect 7882 8630 7986 9487
rect 7851 8588 7986 8630
rect 7886 8501 7986 8588
rect 8064 8500 8212 10479
rect 18237 10713 21805 10747
rect 21895 10713 25463 10747
rect 18175 10318 18209 10654
rect 21833 10318 21867 10654
rect 25491 10318 25525 10654
rect 18237 10225 21805 10259
rect 21895 10225 25463 10259
rect 18175 9830 18209 10166
rect 21833 9830 21867 10166
rect 25491 9830 25525 10166
rect 18237 9737 21805 9771
rect 21895 9737 25463 9771
rect 2688 3829 2862 3875
rect 5629 3873 5741 3875
rect 6371 8356 6562 8370
rect 6371 2963 6473 8356
rect 6473 2963 6507 8356
rect 6507 2963 6562 8356
rect 6731 8215 6907 8249
rect 6647 8019 6681 8187
rect 6957 8019 6991 8187
rect 6731 7957 6907 7991
rect 6647 7761 6681 7929
rect 6957 7761 6991 7929
rect 6731 7699 6907 7733
rect 6647 7503 6681 7671
rect 6957 7503 6991 7671
rect 6731 7441 6907 7475
rect 6647 7245 6681 7413
rect 6957 7245 6991 7413
rect 6731 7183 6907 7217
rect 6647 6987 6681 7155
rect 6957 6987 6991 7155
rect 6731 6925 6907 6959
rect 6647 6729 6681 6897
rect 6957 6729 6991 6897
rect 6731 6667 6907 6701
rect 6647 6471 6681 6639
rect 6957 6471 6991 6639
rect 6731 6409 6907 6443
rect 6647 6213 6681 6381
rect 6957 6213 6991 6381
rect 6731 6151 6907 6185
rect 6647 5955 6681 6123
rect 6957 5955 6991 6123
rect 6731 5893 6907 5927
rect 6647 5697 6681 5865
rect 6957 5697 6991 5865
rect 6731 5635 6907 5669
rect 6647 5439 6681 5607
rect 6957 5439 6991 5607
rect 6731 5377 6907 5411
rect 6647 5181 6681 5349
rect 6957 5181 6991 5349
rect 6731 5119 6907 5153
rect 6647 4923 6681 5091
rect 6957 4923 6991 5091
rect 6731 4861 6907 4895
rect 6647 4665 6681 4833
rect 6957 4665 6991 4833
rect 6731 4603 6907 4637
rect 6647 4407 6681 4575
rect 6957 4407 6991 4575
rect 6731 4345 6907 4379
rect 6647 4149 6681 4317
rect 6957 4149 6991 4317
rect 6731 4087 6907 4121
rect 6647 3891 6681 4059
rect 6957 3891 6991 4059
rect 6731 3829 6907 3863
rect 6647 3633 6681 3801
rect 6957 3633 6991 3801
rect 6731 3571 6907 3605
rect 6647 3375 6681 3543
rect 6957 3375 6991 3543
rect 6731 3313 6907 3347
rect 6647 3117 6681 3285
rect 6957 3117 6991 3285
rect 6731 3055 6907 3089
rect 7518 7899 7694 7933
rect 7425 7503 7459 7871
rect 7753 7503 7787 7871
rect 7518 7441 7694 7475
rect 7518 6609 7694 6643
rect 7425 6213 7459 6581
rect 7753 6213 7787 6581
rect 7518 6151 7694 6185
rect 7518 5319 7694 5353
rect 7425 4923 7459 5291
rect 7753 4923 7787 5291
rect 7518 4861 7694 4895
rect 7518 4029 7694 4063
rect 7425 3633 7459 4001
rect 7753 3633 7787 4001
rect 7518 3571 7694 3605
rect 7518 3448 7694 3482
rect 7425 3052 7459 3420
rect 7753 3052 7787 3420
rect 7518 2990 7694 3024
rect 7965 2945 8104 7940
rect 18058 7235 18634 7269
rect 17974 6239 18008 7207
rect 18684 6239 18718 7207
rect 18058 6177 18634 6211
rect 17832 5573 18385 5667
rect 19447 8832 21815 8866
rect 21905 8832 24273 8866
rect 19385 7606 19419 8782
rect 21843 7606 21877 8782
rect 24301 7606 24335 8782
rect 19447 7522 21815 7556
rect 21905 7522 24273 7556
rect 19446 6957 21814 6991
rect 21904 6957 24272 6991
rect 19384 5731 19418 6907
rect 21842 5731 21876 6907
rect 24300 5731 24334 6907
rect 19446 5647 21814 5681
rect 21904 5647 24272 5681
rect 17834 5343 24768 5432
<< metal1 >>
rect 11788 33012 14404 33018
rect 11788 32803 11800 33012
rect 14392 32809 14404 33012
rect 3389 30890 11211 30896
rect 3389 30801 3401 30890
rect 11199 30801 11211 30890
rect 3389 30795 11211 30801
rect 3519 30533 10966 30539
rect 3519 30499 3728 30533
rect 7296 30499 7386 30533
rect 10954 30499 10966 30533
rect 3519 30493 10966 30499
rect 3519 30440 3719 30493
rect 3519 30104 3666 30440
rect 3700 30104 3719 30440
rect 3519 30091 3719 30104
rect 3519 29060 3605 30091
rect 3896 30051 7135 30493
rect 7318 30440 7364 30452
rect 7304 30104 7314 30440
rect 7368 30104 7378 30440
rect 7318 30092 7364 30104
rect 7558 30051 10797 30493
rect 10962 30440 11164 30453
rect 10962 30104 10982 30440
rect 11016 30104 11164 30440
rect 10962 30093 11164 30104
rect 10976 30092 11022 30093
rect 3716 30045 7308 30051
rect 3716 30011 3728 30045
rect 7296 30011 7308 30045
rect 3716 30005 7308 30011
rect 7374 30045 10966 30051
rect 7374 30011 7386 30045
rect 10954 30011 10966 30045
rect 7374 30005 10966 30011
rect 3633 29952 3719 29964
rect 3633 29921 3666 29952
rect 3700 29921 3719 29952
rect 3709 29616 3719 29921
rect 3633 29603 3719 29616
rect 3896 29563 7135 30005
rect 7318 29952 7364 29964
rect 7304 29616 7314 29952
rect 7368 29616 7378 29952
rect 7318 29604 7364 29616
rect 7558 29563 10797 30005
rect 10964 29952 11050 29964
rect 10964 29911 10982 29952
rect 11016 29911 11050 29952
rect 10964 29616 10974 29911
rect 10964 29563 11050 29616
rect 3716 29557 11050 29563
rect 3716 29523 3728 29557
rect 7296 29523 7386 29557
rect 10954 29523 11050 29557
rect 3716 29517 11050 29523
rect 11078 29245 11164 30093
rect 11790 29401 11800 32803
rect 11965 32803 14404 32809
rect 11965 29401 11975 32803
rect 12188 32609 12560 32615
rect 12188 32575 12200 32609
rect 12548 32575 12560 32609
rect 12188 32569 12560 32575
rect 12626 32609 12998 32615
rect 12626 32575 12638 32609
rect 12986 32575 12998 32609
rect 12626 32569 12998 32575
rect 13064 32609 13436 32615
rect 13064 32575 13076 32609
rect 13424 32575 13436 32609
rect 13064 32569 13436 32575
rect 13502 32609 13874 32615
rect 13502 32575 13514 32609
rect 13862 32575 13874 32609
rect 13502 32569 13874 32575
rect 12132 32516 12178 32528
rect 12132 30540 12138 32516
rect 12172 30540 12178 32516
rect 12112 29540 12122 30540
rect 12186 29540 12196 30540
rect 12132 29528 12178 29540
rect 12260 29490 12465 32569
rect 12570 32516 12616 32528
rect 12547 31916 12557 32516
rect 12629 31916 12639 32516
rect 12570 29540 12576 31916
rect 12610 29540 12616 31916
rect 12570 29528 12616 29540
rect 12713 29490 12918 32569
rect 13008 32516 13054 32528
rect 13008 31777 13014 32516
rect 13048 31777 13054 32516
rect 12989 30777 12999 31777
rect 13063 30777 13073 31777
rect 13008 29540 13014 30777
rect 13048 29540 13054 30777
rect 13008 29528 13054 29540
rect 13149 29490 13354 32569
rect 13446 32516 13492 32528
rect 13423 31916 13433 32516
rect 13505 31916 13515 32516
rect 13446 29540 13452 31916
rect 13486 29540 13492 31916
rect 13446 29528 13492 29540
rect 13589 29490 13794 32569
rect 13884 32516 13930 32528
rect 13884 30540 13890 32516
rect 13924 30540 13930 32516
rect 14174 32230 14328 32242
rect 13865 29540 13875 30540
rect 13939 29540 13949 30540
rect 14174 29750 14180 32230
rect 14322 29750 14328 32230
rect 14174 29738 14328 29750
rect 13884 29528 13930 29540
rect 12190 29487 12200 29490
rect 12188 29441 12200 29487
rect 12480 29487 12490 29490
rect 12628 29487 12638 29490
rect 12480 29481 12560 29487
rect 12548 29447 12560 29481
rect 12190 29438 12200 29441
rect 12480 29441 12560 29447
rect 12626 29441 12638 29487
rect 12918 29487 12928 29490
rect 13066 29487 13076 29490
rect 12918 29481 12998 29487
rect 12986 29447 12998 29481
rect 12480 29438 12490 29441
rect 12628 29438 12638 29441
rect 12918 29441 12998 29447
rect 13064 29441 13076 29487
rect 13356 29487 13366 29490
rect 13504 29487 13514 29490
rect 13356 29481 13436 29487
rect 13424 29447 13436 29481
rect 12918 29438 12928 29441
rect 13066 29438 13076 29441
rect 13356 29441 13436 29447
rect 13502 29441 13514 29487
rect 13794 29487 13804 29490
rect 13794 29481 13874 29487
rect 13862 29447 13874 29481
rect 13356 29438 13366 29441
rect 13504 29438 13514 29441
rect 13794 29441 13874 29447
rect 13794 29438 13804 29441
rect 11794 29389 11971 29401
rect 3633 29238 12200 29245
rect 3942 29230 12200 29238
rect 3942 29163 4441 29230
rect 4790 29227 12200 29230
rect 4790 29163 9505 29227
rect 3942 29160 9505 29163
rect 9854 29160 12200 29227
rect 3942 29154 12200 29160
rect 3633 29145 12200 29154
rect 12300 29145 12886 29245
rect 12986 29145 13324 29245
rect 13424 29145 13514 29245
rect 13614 29145 15339 29245
rect 15621 29145 15631 29245
rect 3519 29044 11060 29060
rect 3519 29040 9925 29044
rect 3519 28973 4868 29040
rect 5217 28977 9925 29040
rect 10274 28977 10639 29044
rect 5217 28974 10639 28977
rect 11029 28974 11060 29044
rect 5217 28973 11060 28974
rect 3519 28960 11060 28973
rect 10974 28936 11060 28960
rect 10974 28836 12448 28936
rect 12548 28836 12638 28936
rect 12738 28836 13076 28936
rect 13176 28836 13762 28936
rect 13862 28836 14019 28936
rect 4926 28652 7318 28658
rect 4926 28618 4938 28652
rect 7306 28618 7318 28652
rect 4926 28612 7318 28618
rect 7384 28652 9776 28658
rect 7384 28618 7396 28652
rect 9764 28618 9776 28652
rect 12258 28638 12268 28641
rect 7384 28612 9776 28618
rect 12188 28632 12268 28638
rect 12548 28638 12558 28641
rect 12696 28638 12706 28641
rect 4870 28568 4916 28580
rect 4822 28000 4832 28568
rect 4918 28000 4928 28568
rect 4822 27434 4876 28000
rect 4870 27392 4876 27434
rect 4910 27434 4928 28000
rect 4910 27392 4916 27434
rect 4870 27380 4916 27392
rect 5574 27354 6659 28612
rect 7328 28568 7374 28580
rect 7328 27743 7334 28568
rect 7368 27743 7374 28568
rect 7316 27424 7326 27743
rect 7378 27424 7388 27743
rect 7328 27392 7334 27424
rect 7368 27392 7374 27424
rect 7328 27380 7374 27392
rect 8078 27354 9165 28612
rect 12188 28598 12200 28632
rect 11811 28583 11971 28595
rect 12188 28592 12268 28598
rect 12258 28589 12268 28592
rect 12548 28592 12560 28638
rect 12626 28632 12706 28638
rect 12986 28638 12996 28641
rect 13134 28638 13144 28641
rect 12626 28598 12638 28632
rect 12626 28592 12706 28598
rect 12548 28589 12558 28592
rect 12696 28589 12706 28592
rect 12986 28592 12998 28638
rect 13064 28632 13144 28638
rect 13424 28638 13434 28641
rect 13572 28638 13582 28641
rect 13064 28598 13076 28632
rect 13064 28592 13144 28598
rect 12986 28589 12996 28592
rect 13134 28589 13144 28592
rect 13424 28592 13436 28638
rect 13502 28632 13582 28638
rect 13862 28638 13872 28641
rect 13502 28598 13514 28632
rect 13502 28592 13582 28598
rect 13424 28589 13434 28592
rect 13572 28589 13582 28592
rect 13862 28592 13874 28638
rect 13862 28589 13872 28592
rect 9786 28568 9832 28580
rect 9774 28000 9784 28568
rect 9870 28000 9880 28568
rect 9774 27447 9792 28000
rect 9786 27392 9792 27447
rect 9826 27447 9880 28000
rect 9826 27392 9832 27447
rect 9786 27380 9832 27392
rect 4932 27348 4942 27354
rect 4926 27342 4942 27348
rect 5152 27348 7316 27354
rect 7386 27348 9554 27354
rect 5152 27342 7318 27348
rect 4926 27308 4938 27342
rect 7306 27308 7318 27342
rect 4926 27302 4942 27308
rect 4932 27297 4942 27302
rect 5152 27302 7318 27308
rect 7384 27342 9554 27348
rect 9764 27348 9774 27354
rect 7384 27308 7396 27342
rect 7384 27302 9554 27308
rect 5152 27297 7316 27302
rect 7386 27297 9554 27302
rect 9764 27302 9776 27348
rect 9764 27297 9774 27302
rect 4942 27236 7395 27240
rect 4942 27179 4965 27236
rect 5152 27179 7395 27236
rect 4942 27176 7395 27179
rect 7596 27176 7605 27240
rect 4942 27161 7605 27176
rect 3539 27061 3549 27072
rect 3537 27017 3549 27061
rect 4125 27061 4135 27072
rect 4125 27017 4137 27061
rect 3537 27015 4137 27017
rect 3459 26993 3505 27005
rect 3459 26025 3465 26993
rect 3499 26806 3505 26993
rect 4169 26993 4228 27005
rect 4169 26824 4175 26993
rect 4209 26824 4228 26993
rect 7095 26923 9764 26943
rect 7095 26921 9554 26923
rect 7305 26866 9554 26921
rect 7305 26864 9764 26866
rect 7095 26854 9764 26864
rect 4157 26806 4167 26824
rect 3499 26209 4167 26806
rect 3499 26025 3505 26209
rect 4157 26025 4167 26209
rect 4219 26025 4229 26824
rect 4927 26783 7095 26789
rect 4925 26777 7095 26783
rect 7305 26783 7315 26789
rect 7385 26783 7395 26788
rect 4925 26743 4937 26777
rect 4925 26737 7095 26743
rect 4927 26732 7095 26737
rect 7305 26737 7317 26783
rect 7383 26737 7395 26783
rect 7605 26783 9773 26788
rect 7605 26777 9775 26783
rect 9763 26743 9775 26777
rect 7305 26732 7315 26737
rect 4869 26693 4915 26705
rect 3459 26013 3505 26025
rect 4169 26013 4228 26025
rect 3537 25997 4137 26003
rect 3537 25963 3549 25997
rect 4125 25963 4137 25997
rect 3537 25957 4137 25963
rect 4716 25621 4765 26693
rect 4917 25621 4927 26693
rect 4716 25552 4875 25621
rect 4869 25517 4875 25552
rect 4909 25552 4927 25621
rect 4909 25517 4915 25552
rect 4869 25505 4915 25517
rect 5569 25474 6656 26732
rect 7385 26731 7395 26737
rect 7605 26737 9775 26743
rect 7605 26731 9773 26737
rect 7327 26693 7373 26705
rect 7327 26662 7333 26693
rect 7367 26662 7373 26693
rect 7315 26343 7325 26662
rect 7377 26343 7387 26662
rect 7327 25517 7333 26343
rect 7367 25517 7373 26343
rect 7327 25505 7373 25517
rect 3311 25453 3888 25459
rect 3311 25359 3323 25453
rect 3876 25359 3888 25453
rect 4925 25422 4937 25474
rect 5417 25467 7317 25474
rect 7385 25473 7395 25475
rect 7305 25433 7317 25467
rect 5417 25422 7317 25433
rect 7383 25427 7395 25473
rect 7875 25473 7885 25475
rect 8069 25473 9156 26731
rect 9785 26693 9831 26705
rect 9772 25621 9782 26693
rect 9934 25621 9944 26693
rect 9785 25517 9791 25621
rect 9825 25517 9831 25621
rect 9785 25505 9831 25517
rect 7875 25467 9775 25473
rect 9763 25433 9775 25467
rect 7385 25423 7395 25427
rect 7875 25427 9775 25433
rect 7875 25423 7885 25427
rect 11807 25407 11817 28583
rect 3311 25353 3888 25359
rect 11806 25231 11816 25407
rect 11965 25380 11975 28583
rect 12132 28539 12178 28551
rect 12113 27539 12123 28539
rect 12187 27539 12197 28539
rect 12132 25563 12138 27539
rect 12172 25563 12178 27539
rect 12132 25551 12178 25563
rect 12264 25510 12469 28589
rect 12570 28539 12616 28551
rect 12570 26163 12576 28539
rect 12610 26163 12616 28539
rect 12547 25563 12557 26163
rect 12629 25563 12639 26163
rect 12570 25551 12616 25563
rect 12717 25510 12922 28589
rect 13008 28539 13054 28551
rect 13008 27379 13014 28539
rect 13048 27379 13054 28539
rect 12989 26379 12999 27379
rect 13063 26379 13073 27379
rect 13008 25563 13014 26379
rect 13048 25563 13054 26379
rect 13008 25551 13054 25563
rect 13153 25510 13358 28589
rect 13446 28539 13492 28551
rect 13446 26163 13452 28539
rect 13486 26163 13492 28539
rect 13422 25563 13432 26163
rect 13504 25563 13514 26163
rect 13446 25551 13492 25563
rect 13585 25510 13790 28589
rect 13884 28539 13930 28551
rect 13865 27539 13875 28539
rect 13939 27539 13949 28539
rect 25397 28163 25668 28170
rect 20688 28158 25668 28163
rect 20688 28157 25403 28158
rect 14190 27997 14344 28009
rect 13884 25563 13890 27539
rect 13924 25563 13930 27539
rect 13884 25551 13930 25563
rect 14190 25517 14196 27997
rect 14338 27505 14344 27997
rect 20688 27792 20700 28157
rect 25662 27793 25672 28158
rect 25504 27792 25546 27793
rect 20688 27786 20762 27792
rect 18845 27505 19144 27510
rect 14338 27499 19144 27505
rect 19128 27498 19144 27499
rect 14338 27201 16600 27207
rect 14338 25517 14344 27201
rect 12188 25504 12560 25510
rect 12188 25470 12200 25504
rect 12548 25470 12560 25504
rect 12188 25464 12560 25470
rect 12626 25504 12998 25510
rect 12626 25470 12638 25504
rect 12986 25470 12998 25504
rect 12626 25464 12998 25470
rect 13064 25504 13436 25510
rect 13064 25470 13076 25504
rect 13424 25470 13436 25504
rect 13064 25464 13436 25470
rect 13502 25504 13874 25510
rect 14190 25505 14344 25517
rect 13502 25470 13514 25504
rect 13862 25470 13874 25504
rect 13502 25464 13874 25470
rect 11965 25374 14393 25380
rect 11810 25230 11929 25231
rect 14381 25230 14393 25374
rect 11810 25224 14393 25230
rect 3313 25218 10271 25224
rect 11810 25219 11971 25224
rect 3313 25129 3325 25218
rect 10259 25129 10271 25218
rect 16594 25217 16600 27201
rect 16833 27201 18851 27207
rect 16833 25457 16839 27201
rect 17017 27078 17369 27084
rect 17017 27044 17029 27078
rect 17357 27044 17369 27078
rect 17017 27038 17369 27044
rect 17435 27078 17787 27084
rect 17435 27044 17447 27078
rect 17775 27044 17787 27078
rect 17435 27038 17787 27044
rect 17853 27078 18205 27084
rect 17853 27044 17865 27078
rect 18193 27044 18205 27078
rect 17853 27038 18205 27044
rect 18271 27078 18623 27084
rect 18271 27044 18283 27078
rect 18611 27044 18623 27078
rect 18271 27038 18623 27044
rect 16961 26985 17007 26997
rect 16948 25985 16958 26985
rect 17010 25985 17020 26985
rect 16961 25609 16967 25985
rect 17001 25609 17007 25985
rect 16961 25597 17007 25609
rect 17085 25556 17286 27038
rect 17379 26985 17425 26997
rect 17379 26609 17385 26985
rect 17419 26609 17425 26985
rect 17366 25609 17376 26609
rect 17428 25609 17438 26609
rect 17379 25597 17425 25609
rect 17504 25556 17705 27038
rect 17797 26985 17843 26997
rect 17784 25985 17794 26985
rect 17846 25985 17856 26985
rect 17797 25609 17803 25985
rect 17837 25609 17843 25985
rect 17797 25597 17843 25609
rect 17927 25556 18128 27038
rect 18215 26985 18261 26997
rect 18215 26609 18221 26985
rect 18255 26609 18261 26985
rect 18202 25609 18212 26609
rect 18264 25609 18274 26609
rect 18215 25597 18261 25609
rect 18333 25556 18534 27038
rect 18633 26985 18679 26997
rect 18620 25985 18630 26985
rect 18682 25985 18692 26985
rect 18633 25609 18639 25985
rect 18673 25609 18679 25985
rect 18841 25691 18851 27201
rect 19138 25691 19148 27498
rect 18845 25679 19144 25691
rect 18633 25597 18679 25609
rect 18828 25556 18838 25565
rect 17017 25550 18838 25556
rect 17017 25516 17029 25550
rect 17357 25516 17447 25550
rect 17775 25516 17865 25550
rect 18193 25516 18283 25550
rect 18611 25516 18838 25550
rect 17017 25510 18838 25516
rect 18828 25506 18838 25510
rect 18962 25506 18972 25565
rect 20752 25500 20762 27786
rect 20879 27786 25546 27792
rect 20879 25596 20889 27786
rect 25397 27781 25546 27786
rect 21054 27623 22102 27629
rect 21054 27589 21122 27623
rect 22090 27589 22102 27623
rect 21054 27583 22102 27589
rect 22168 27623 24218 27629
rect 22168 27589 22180 27623
rect 23148 27589 23238 27623
rect 24206 27589 24218 27623
rect 22168 27583 24218 27589
rect 24284 27623 25332 27629
rect 24284 27589 24296 27623
rect 25264 27589 25332 27623
rect 24284 27583 25332 27589
rect 21054 27530 21100 27583
rect 21054 27254 21060 27530
rect 21094 27254 21100 27530
rect 21035 27054 21045 27254
rect 21109 27054 21119 27254
rect 21054 27001 21100 27054
rect 21255 27004 21908 27583
rect 22112 27530 22158 27542
rect 22099 27230 22109 27530
rect 22161 27230 22171 27530
rect 22112 27054 22118 27230
rect 22152 27054 22158 27230
rect 22112 27042 22158 27054
rect 22341 27004 22994 27583
rect 23170 27530 23216 27583
rect 23151 27330 23161 27530
rect 23225 27330 23235 27530
rect 23170 27054 23176 27330
rect 23210 27054 23216 27330
rect 23170 27004 23216 27054
rect 23411 27005 24064 27583
rect 24228 27530 24274 27542
rect 24215 27230 24225 27530
rect 24277 27230 24287 27530
rect 24228 27054 24234 27230
rect 24268 27054 24274 27230
rect 24228 27042 24274 27054
rect 21255 27001 21450 27004
rect 21054 26995 21450 27001
rect 22090 27001 22100 27004
rect 22341 27001 22508 27004
rect 21054 26961 21122 26995
rect 21054 26955 21450 26961
rect 21440 26952 21450 26955
rect 22090 26955 22102 27001
rect 22168 26995 22508 27001
rect 23148 27001 23231 27004
rect 23411 27001 23566 27005
rect 23148 26995 23566 27001
rect 24206 27001 24216 27005
rect 24444 27004 25097 27583
rect 25286 27530 25332 27583
rect 25286 27254 25292 27530
rect 25326 27254 25332 27530
rect 25267 27054 25277 27254
rect 25341 27054 25351 27254
rect 25286 27042 25332 27054
rect 24444 27001 24624 27004
rect 22168 26961 22180 26995
rect 23148 26961 23238 26995
rect 22168 26955 22508 26961
rect 22090 26952 22100 26955
rect 22498 26952 22508 26955
rect 23148 26955 23566 26961
rect 23148 26952 23231 26955
rect 23556 26953 23566 26955
rect 24206 26955 24218 27001
rect 24284 26995 24624 27001
rect 25264 27001 25274 27004
rect 24284 26961 24296 26995
rect 24284 26955 24624 26961
rect 24206 26953 24216 26955
rect 24614 26952 24624 26955
rect 25264 26955 25276 27001
rect 25536 26979 25546 27781
rect 25643 27781 25668 27793
rect 25643 26979 25653 27781
rect 25540 26967 25649 26979
rect 25264 26952 25274 26955
rect 21103 26756 21990 26856
rect 22090 26756 22180 26856
rect 22280 26756 23238 26856
rect 23338 26756 25164 26856
rect 25264 26756 25879 26856
rect 21106 26574 21122 26674
rect 21222 26574 23048 26674
rect 23148 26574 24106 26674
rect 24206 26574 24296 26674
rect 24396 26574 25524 26674
rect 21054 26470 21100 26471
rect 21054 26418 21122 26470
rect 21762 26467 21772 26470
rect 22170 26467 22180 26470
rect 21762 26461 22102 26467
rect 22090 26427 22102 26461
rect 21762 26421 22102 26427
rect 22168 26421 22180 26467
rect 22820 26467 22830 26470
rect 23228 26467 23238 26470
rect 22820 26461 23238 26467
rect 23878 26467 23888 26470
rect 24286 26467 24296 26470
rect 23878 26461 24218 26467
rect 23148 26427 23238 26461
rect 24206 26427 24218 26461
rect 21762 26418 21945 26421
rect 22170 26418 22180 26421
rect 22820 26421 23238 26427
rect 22820 26418 22977 26421
rect 21054 26417 21132 26418
rect 21054 26368 21100 26417
rect 21035 26168 21045 26368
rect 21109 26168 21119 26368
rect 21054 25892 21060 26168
rect 21094 25892 21100 26168
rect 21054 25839 21100 25892
rect 21292 25839 21945 26418
rect 22112 26368 22158 26380
rect 22112 26192 22118 26368
rect 22152 26192 22158 26368
rect 22099 25892 22109 26192
rect 22161 25892 22171 26192
rect 22112 25880 22158 25892
rect 22324 25839 22977 26418
rect 23170 26418 23238 26421
rect 23878 26421 24218 26427
rect 24284 26421 24296 26467
rect 24936 26467 24946 26470
rect 24936 26461 25332 26467
rect 25264 26427 25332 26461
rect 23878 26418 24088 26421
rect 24286 26418 24296 26421
rect 24936 26421 25332 26427
rect 24936 26418 25126 26421
rect 23170 26368 23216 26418
rect 23170 26092 23176 26368
rect 23210 26092 23216 26368
rect 23151 25892 23161 26092
rect 23225 25892 23235 26092
rect 23170 25839 23216 25892
rect 23435 25839 24088 26418
rect 24228 26368 24274 26380
rect 24228 26192 24234 26368
rect 24268 26192 24274 26368
rect 24215 25892 24225 26192
rect 24277 25892 24287 26192
rect 24228 25880 24274 25892
rect 24473 25839 25126 26418
rect 25286 26368 25332 26421
rect 25267 26168 25277 26368
rect 25341 26168 25351 26368
rect 25286 25892 25292 26168
rect 25326 25892 25332 26168
rect 25286 25839 25332 25892
rect 21054 25833 22102 25839
rect 21054 25799 21122 25833
rect 22090 25799 22102 25833
rect 21054 25793 22102 25799
rect 22168 25833 24218 25839
rect 22168 25799 22180 25833
rect 23148 25799 23238 25833
rect 24206 25799 24218 25833
rect 22168 25793 24218 25799
rect 24284 25833 25332 25839
rect 24284 25799 24296 25833
rect 25264 25799 25332 25833
rect 24284 25793 25332 25799
rect 20879 25590 25323 25596
rect 20756 25493 20797 25500
rect 20756 25488 25207 25493
rect 20785 25487 25207 25488
rect 16833 25451 18760 25457
rect 16594 25215 16685 25217
rect 18748 25215 18760 25451
rect 22114 25366 22184 25372
rect 24187 25366 24275 25372
rect 22114 25360 24275 25366
rect 16594 25209 18760 25215
rect 16594 25205 16839 25209
rect 3313 25123 10271 25129
rect 19692 24929 19820 24948
rect 11866 24892 12025 24904
rect 11862 23596 11872 24892
rect 12019 24890 12029 24892
rect 12019 24889 12160 24890
rect 19682 24889 19692 24929
rect 12019 24884 19692 24889
rect 12148 24883 19692 24884
rect 11860 23392 11872 23596
rect 12019 24774 19692 24780
rect 12019 23596 12029 24774
rect 19682 24746 19692 24774
rect 19839 24746 19849 24929
rect 22110 24719 22120 25360
rect 22178 25251 24193 25257
rect 22178 24719 22188 25251
rect 22295 25167 22687 25173
rect 22295 25133 22307 25167
rect 22675 25133 22687 25167
rect 22295 25127 22687 25133
rect 22753 25167 23145 25173
rect 22753 25133 22765 25167
rect 23133 25133 23145 25167
rect 22753 25127 23145 25133
rect 23211 25167 23603 25173
rect 23211 25133 23223 25167
rect 23591 25133 23603 25167
rect 23211 25127 23603 25133
rect 23669 25167 24061 25173
rect 23669 25133 23681 25167
rect 24049 25133 24061 25167
rect 23669 25127 24061 25133
rect 22239 25083 22285 25095
rect 22114 24707 22184 24719
rect 22239 24654 22245 25083
rect 22279 24654 22285 25083
rect 12198 24597 14070 24603
rect 12198 24563 12210 24597
rect 14058 24563 14070 24597
rect 12198 24557 14070 24563
rect 14136 24597 17946 24603
rect 14136 24563 14148 24597
rect 15996 24563 16086 24597
rect 17934 24563 17946 24597
rect 14136 24557 17946 24563
rect 18012 24597 19884 24603
rect 18012 24563 18024 24597
rect 19872 24563 19884 24597
rect 18012 24557 19884 24563
rect 12142 24513 12188 24525
rect 12123 24413 12133 24513
rect 12197 24413 12207 24513
rect 12142 24237 12148 24413
rect 12182 24237 12188 24413
rect 12142 24225 12188 24237
rect 12418 24193 13837 24557
rect 14080 24513 14126 24525
rect 14067 24413 14077 24513
rect 14129 24413 14139 24513
rect 14080 24237 14086 24413
rect 14120 24237 14126 24413
rect 14080 24225 14126 24237
rect 14452 24193 15871 24557
rect 16018 24513 16064 24557
rect 16018 24337 16024 24513
rect 16058 24337 16064 24513
rect 15999 24237 16009 24337
rect 16073 24237 16083 24337
rect 16018 24225 16064 24237
rect 16281 24193 17700 24557
rect 17956 24513 18002 24525
rect 17943 24413 17953 24513
rect 18005 24413 18015 24513
rect 17956 24237 17962 24413
rect 17996 24237 18002 24413
rect 17956 24225 18002 24237
rect 18251 24193 19670 24557
rect 19894 24513 19940 24525
rect 22203 24517 22213 24654
rect 22307 24517 22317 24654
rect 19875 24413 19885 24513
rect 19949 24413 19959 24513
rect 22239 24507 22245 24517
rect 22279 24507 22285 24517
rect 22239 24495 22285 24507
rect 22371 24466 22592 25127
rect 22697 25083 22743 25095
rect 22684 24923 22694 25083
rect 22746 24923 22756 25083
rect 22697 24507 22703 24923
rect 22737 24507 22743 24923
rect 22697 24495 22743 24507
rect 22830 24466 23051 25127
rect 23155 25083 23201 25095
rect 23155 24912 23161 25083
rect 23195 24912 23201 25083
rect 23122 24775 23132 24912
rect 23226 24775 23236 24912
rect 23155 24507 23161 24775
rect 23195 24507 23201 24775
rect 23155 24495 23201 24507
rect 23293 24466 23514 25127
rect 23613 25083 23659 25095
rect 23600 24923 23610 25083
rect 23662 24923 23672 25083
rect 23613 24507 23619 24923
rect 23653 24507 23659 24923
rect 23613 24495 23659 24507
rect 23747 24466 23968 25127
rect 24071 25083 24117 25095
rect 24071 24654 24077 25083
rect 24111 24654 24117 25083
rect 24038 24517 24048 24654
rect 24142 24517 24152 24654
rect 24071 24507 24077 24517
rect 24111 24507 24117 24517
rect 24071 24495 24117 24507
rect 22371 24463 22475 24466
rect 22295 24457 22475 24463
rect 22675 24463 22685 24466
rect 22830 24463 22933 24466
rect 22295 24423 22307 24457
rect 22295 24417 22475 24423
rect 22465 24414 22475 24417
rect 22675 24417 22687 24463
rect 22753 24457 22933 24463
rect 23133 24463 23143 24466
rect 23293 24463 23391 24466
rect 22753 24423 22765 24457
rect 22753 24417 22933 24423
rect 22675 24414 22685 24417
rect 22923 24414 22933 24417
rect 23133 24417 23145 24463
rect 23211 24457 23391 24463
rect 23591 24463 23601 24466
rect 23747 24463 23849 24466
rect 23211 24423 23223 24457
rect 23211 24417 23391 24423
rect 23133 24414 23143 24417
rect 23381 24414 23391 24417
rect 23591 24417 23603 24463
rect 23669 24457 23849 24463
rect 24049 24463 24059 24466
rect 23669 24423 23681 24457
rect 23669 24417 23849 24423
rect 23591 24414 23601 24417
rect 23839 24414 23849 24417
rect 24049 24417 24061 24463
rect 24049 24414 24059 24417
rect 19894 24237 19900 24413
rect 19934 24237 19940 24413
rect 20726 24242 20736 24342
rect 20819 24242 22575 24342
rect 22675 24242 22765 24342
rect 22865 24242 23223 24342
rect 23323 24242 23949 24342
rect 24049 24242 24094 24342
rect 19894 24225 19940 24237
rect 12198 24187 19884 24193
rect 12198 24153 12210 24187
rect 14058 24153 14148 24187
rect 15996 24153 16086 24187
rect 17934 24153 18024 24187
rect 19872 24153 19884 24187
rect 12198 24147 19884 24153
rect 12142 24103 12188 24115
rect 12142 23927 12148 24103
rect 12182 23927 12188 24103
rect 12123 23827 12133 23927
rect 12197 23827 12207 23927
rect 12142 23783 12188 23827
rect 12422 23783 13841 24147
rect 14080 24103 14126 24115
rect 14080 23927 14086 24103
rect 14120 23927 14126 24103
rect 14067 23827 14077 23927
rect 14129 23827 14139 23927
rect 14080 23815 14126 23827
rect 14448 23783 15867 24147
rect 16018 24103 16064 24115
rect 15999 24003 16009 24103
rect 16073 24003 16083 24103
rect 16018 23827 16024 24003
rect 16058 23827 16064 24003
rect 16018 23815 16064 23827
rect 16281 23783 17700 24147
rect 17956 24103 18002 24115
rect 17956 23927 17962 24103
rect 17996 23927 18002 24103
rect 17943 23827 17953 23927
rect 18005 23827 18015 23927
rect 17956 23815 18002 23827
rect 18251 23783 19670 24147
rect 19894 24103 19940 24115
rect 19894 23927 19900 24103
rect 19934 23927 19940 24103
rect 20716 24056 20726 24156
rect 20839 24056 22307 24156
rect 22407 24056 23033 24156
rect 23133 24056 23491 24156
rect 23591 24056 23681 24156
rect 23781 24056 24094 24156
rect 22297 23966 22307 23969
rect 19875 23827 19885 23927
rect 19949 23827 19959 23927
rect 22295 23920 22307 23966
rect 22507 23966 22517 23969
rect 22755 23966 22765 23969
rect 22507 23960 22687 23966
rect 22675 23926 22687 23960
rect 22297 23917 22307 23920
rect 22507 23920 22687 23926
rect 22753 23920 22765 23966
rect 22965 23966 22975 23969
rect 23213 23966 23223 23969
rect 22965 23960 23145 23966
rect 23133 23926 23145 23960
rect 22507 23917 22594 23920
rect 22755 23917 22765 23920
rect 22965 23920 23145 23926
rect 23211 23920 23223 23966
rect 23423 23966 23433 23969
rect 23671 23966 23681 23969
rect 23423 23960 23603 23966
rect 23591 23926 23603 23960
rect 22965 23917 23057 23920
rect 23213 23917 23223 23920
rect 23423 23920 23603 23926
rect 23669 23920 23681 23966
rect 23881 23966 23891 23969
rect 23881 23960 24061 23966
rect 24049 23926 24061 23960
rect 23423 23917 23502 23920
rect 23671 23917 23681 23920
rect 23881 23920 24061 23926
rect 23881 23917 23972 23920
rect 22239 23876 22285 23888
rect 22239 23865 22245 23876
rect 22279 23865 22285 23876
rect 19894 23783 19940 23827
rect 12142 23777 14070 23783
rect 12142 23743 12210 23777
rect 14058 23743 14070 23777
rect 12142 23737 14070 23743
rect 14136 23777 16008 23783
rect 14136 23743 14148 23777
rect 15996 23743 16008 23777
rect 14136 23737 16008 23743
rect 16074 23777 17946 23783
rect 16074 23743 16086 23777
rect 17934 23743 17946 23777
rect 16074 23737 17946 23743
rect 18012 23777 19940 23783
rect 18012 23743 18024 23777
rect 19872 23743 19940 23777
rect 18012 23737 19940 23743
rect 22204 23728 22214 23865
rect 22308 23728 22318 23865
rect 22105 23683 22191 23695
rect 12019 23595 12125 23596
rect 12019 23590 19803 23595
rect 12113 23589 19803 23590
rect 19791 23392 19803 23589
rect 11860 23386 19803 23392
rect 22101 23064 22111 23683
rect 22060 23052 22111 23064
rect 22185 23064 22195 23683
rect 22239 23300 22245 23728
rect 22279 23300 22285 23728
rect 22239 23288 22285 23300
rect 22373 23256 22594 23917
rect 22697 23876 22743 23888
rect 22697 23460 22703 23876
rect 22737 23460 22743 23876
rect 22684 23300 22694 23460
rect 22746 23300 22756 23460
rect 22697 23288 22743 23300
rect 22836 23256 23057 23917
rect 23155 23876 23201 23888
rect 23155 23654 23161 23876
rect 23195 23654 23201 23876
rect 23121 23517 23131 23654
rect 23225 23517 23235 23654
rect 23155 23300 23161 23517
rect 23195 23300 23201 23517
rect 23155 23288 23201 23300
rect 23281 23256 23502 23917
rect 23613 23876 23659 23888
rect 23613 23460 23619 23876
rect 23653 23460 23659 23876
rect 23600 23300 23610 23460
rect 23662 23300 23672 23460
rect 23613 23288 23659 23300
rect 23751 23256 23972 23917
rect 24071 23876 24117 23888
rect 24071 23865 24077 23876
rect 24111 23865 24117 23876
rect 24036 23728 24046 23865
rect 24140 23728 24150 23865
rect 24071 23300 24077 23728
rect 24111 23300 24117 23728
rect 24071 23288 24117 23300
rect 22295 23250 22687 23256
rect 22295 23216 22307 23250
rect 22675 23216 22687 23250
rect 22295 23210 22687 23216
rect 22753 23250 23145 23256
rect 22753 23216 22765 23250
rect 23133 23216 23145 23250
rect 22753 23210 23145 23216
rect 23211 23250 23603 23256
rect 23211 23216 23223 23250
rect 23591 23216 23603 23250
rect 23211 23210 23603 23216
rect 23669 23250 24061 23256
rect 23669 23216 23681 23250
rect 24049 23216 24061 23250
rect 23669 23210 24061 23216
rect 22185 23058 22299 23064
rect 24187 23058 24193 25251
rect 22185 23052 24193 23058
rect 24269 23058 24275 25360
rect 25197 24334 25207 25487
rect 25311 25487 25323 25590
rect 25311 24334 25321 25487
rect 25424 25058 25524 26574
rect 25424 25024 25455 25058
rect 25493 25024 25524 25058
rect 25424 25018 25524 25024
rect 25779 25058 25879 26756
rect 25779 25024 25811 25058
rect 25849 25024 25879 25058
rect 25779 25018 25879 25024
rect 25387 24965 25433 24977
rect 25515 24965 25561 24977
rect 25743 24965 25789 24977
rect 25871 24965 25917 24977
rect 25374 24765 25384 24965
rect 25436 24765 25446 24965
rect 25387 24469 25393 24765
rect 25427 24469 25433 24765
rect 25515 24669 25521 24965
rect 25555 24669 25561 24965
rect 25730 24765 25740 24965
rect 25792 24765 25802 24965
rect 25502 24469 25512 24669
rect 25564 24469 25574 24669
rect 25743 24469 25749 24765
rect 25783 24469 25789 24765
rect 25871 24669 25877 24965
rect 25911 24669 25917 24965
rect 25858 24469 25868 24669
rect 25920 24469 25930 24669
rect 25387 24457 25433 24469
rect 25515 24457 25561 24469
rect 25743 24457 25789 24469
rect 25871 24457 25917 24469
rect 25441 24410 25506 24417
rect 25441 24376 25455 24410
rect 25493 24376 25506 24410
rect 25441 24359 25506 24376
rect 25799 24410 25861 24416
rect 25799 24376 25811 24410
rect 25849 24376 25861 24410
rect 25799 24345 25861 24376
rect 25201 24322 25317 24334
rect 25502 24050 25512 24083
rect 25465 24044 25512 24050
rect 25465 24010 25477 24044
rect 25511 24010 25512 24044
rect 25465 24004 25512 24010
rect 25564 24050 25574 24083
rect 25564 24044 25879 24050
rect 25564 24010 25833 24044
rect 25867 24010 25879 24044
rect 25564 24004 25879 24010
rect 25521 23972 25555 24004
rect 25427 23960 25473 23972
rect 25427 23855 25433 23960
rect 25467 23855 25473 23960
rect 25515 23960 25561 23972
rect 25414 23784 25424 23855
rect 25476 23784 25486 23855
rect 25515 23784 25521 23960
rect 25555 23784 25561 23960
rect 25783 23960 25829 23972
rect 25871 23960 25917 23972
rect 25783 23855 25789 23960
rect 25823 23855 25829 23960
rect 25858 23889 25868 23960
rect 25920 23889 25930 23960
rect 25770 23784 25780 23855
rect 25832 23784 25842 23855
rect 25871 23784 25877 23889
rect 25911 23784 25917 23889
rect 25427 23772 25473 23784
rect 25515 23772 25561 23784
rect 25783 23772 25829 23784
rect 25871 23772 25917 23784
rect 25465 23734 25879 23740
rect 25465 23700 25477 23734
rect 25511 23700 25833 23734
rect 25867 23700 25879 23734
rect 25465 23694 25879 23700
rect 24599 23500 26001 23506
rect 24599 23222 24611 23500
rect 25989 23228 26001 23500
rect 24605 23064 24611 23222
rect 24536 23058 24611 23064
rect 24269 23052 24611 23058
rect 24731 23222 26001 23228
rect 17324 22497 17475 22507
rect 15730 22467 15933 22479
rect 12047 21700 12233 21712
rect 12047 15122 12053 21700
rect 12227 15122 12233 21700
rect 14988 21656 15112 21668
rect 12478 21585 12678 21595
rect 12466 21530 12478 21576
rect 14535 21579 14735 21589
rect 12678 21570 13266 21576
rect 13254 21536 13266 21570
rect 13947 21570 14535 21576
rect 12678 21530 13266 21536
rect 13521 21556 13573 21566
rect 12388 21508 12434 21520
rect 12478 21511 12678 21521
rect 13298 21518 13344 21520
rect 12388 21340 12394 21508
rect 12428 21469 12434 21508
rect 13295 21508 13347 21518
rect 12428 21408 13295 21469
rect 12428 21381 13304 21408
rect 12428 21340 12434 21381
rect 12388 21250 12434 21340
rect 13298 21340 13304 21381
rect 13338 21398 13347 21408
rect 13338 21340 13344 21398
rect 13054 21323 13254 21333
rect 12466 21312 13054 21318
rect 12466 21278 12478 21312
rect 12466 21272 13054 21278
rect 13254 21272 13266 21318
rect 13054 21257 13254 21267
rect 12388 21082 12394 21250
rect 12428 21226 12434 21250
rect 13298 21250 13344 21340
rect 13298 21226 13304 21250
rect 12428 21138 13304 21226
rect 12428 21082 12434 21138
rect 12388 21070 12434 21082
rect 13298 21082 13304 21138
rect 13338 21082 13344 21250
rect 12830 21063 12930 21073
rect 13298 21070 13344 21082
rect 13521 21298 13573 21456
rect 12466 21054 12830 21060
rect 12930 21054 13266 21060
rect 12466 21020 12478 21054
rect 13254 21020 13266 21054
rect 12466 21014 12830 21020
rect 12930 21014 13266 21020
rect 12388 20992 12434 21004
rect 12830 21001 12930 21011
rect 13298 21002 13344 21004
rect 12388 20824 12394 20992
rect 12428 20952 12434 20992
rect 13295 20992 13347 21002
rect 12428 20934 13295 20952
rect 12428 20882 12824 20934
rect 12929 20892 13295 20934
rect 12929 20882 13304 20892
rect 12428 20864 13304 20882
rect 12428 20824 12434 20864
rect 12388 20734 12434 20824
rect 13298 20824 13304 20864
rect 13338 20882 13347 20892
rect 13338 20824 13344 20882
rect 12478 20805 12678 20815
rect 12466 20756 12478 20802
rect 12678 20796 13266 20802
rect 13254 20762 13266 20796
rect 12678 20756 13266 20762
rect 12478 20743 12678 20753
rect 12388 20566 12394 20734
rect 12428 20695 12434 20734
rect 13298 20734 13344 20824
rect 13298 20695 13304 20734
rect 12428 20672 13304 20695
rect 12428 20620 12827 20672
rect 12927 20620 13304 20672
rect 12428 20607 13304 20620
rect 12428 20566 12434 20607
rect 12388 20554 12434 20566
rect 13298 20566 13304 20607
rect 13338 20566 13344 20734
rect 12830 20547 12930 20557
rect 13298 20554 13344 20566
rect 12466 20538 12830 20544
rect 12930 20538 13266 20544
rect 12466 20504 12478 20538
rect 13254 20504 13266 20538
rect 12466 20498 12830 20504
rect 12930 20498 13266 20504
rect 13521 20524 13573 21198
rect 12388 20476 12434 20488
rect 12830 20485 12930 20495
rect 13298 20486 13344 20488
rect 12388 20308 12394 20476
rect 12428 20429 12434 20476
rect 13295 20476 13347 20486
rect 12428 20351 13295 20429
rect 12428 20341 13304 20351
rect 12428 20308 12434 20341
rect 12388 20218 12434 20308
rect 13298 20308 13304 20341
rect 13338 20345 13347 20351
rect 13338 20308 13344 20345
rect 13054 20291 13254 20301
rect 12466 20280 13054 20286
rect 12466 20246 12478 20280
rect 12466 20240 13054 20246
rect 13254 20240 13266 20286
rect 13054 20225 13254 20235
rect 12388 20050 12394 20218
rect 12428 20178 12434 20218
rect 13298 20218 13344 20308
rect 13298 20178 13304 20218
rect 12428 20090 13304 20178
rect 12428 20050 12434 20090
rect 12388 19960 12434 20050
rect 13298 20050 13304 20090
rect 13338 20050 13344 20218
rect 12478 20037 12678 20047
rect 12466 19982 12478 20028
rect 12678 20022 13266 20028
rect 13254 19988 13266 20022
rect 12678 19982 13266 19988
rect 12478 19963 12678 19973
rect 12388 19792 12394 19960
rect 12428 19913 12434 19960
rect 13298 19960 13344 20050
rect 13298 19913 13304 19960
rect 12428 19825 13304 19913
rect 12428 19792 12434 19825
rect 12388 19702 12434 19792
rect 13298 19792 13304 19825
rect 13338 19792 13344 19960
rect 13054 19775 13254 19785
rect 12466 19764 13054 19770
rect 12466 19730 12478 19764
rect 12466 19724 13054 19730
rect 13254 19724 13266 19770
rect 13054 19709 13254 19719
rect 12388 19534 12394 19702
rect 12428 19669 12434 19702
rect 13298 19702 13344 19792
rect 13298 19669 13304 19702
rect 12428 19581 13304 19669
rect 12428 19534 12434 19581
rect 12388 19522 12434 19534
rect 13298 19534 13304 19581
rect 13338 19534 13344 19702
rect 12830 19515 12930 19525
rect 13298 19522 13344 19534
rect 13521 19750 13573 20424
rect 12466 19506 12830 19512
rect 12930 19506 13266 19512
rect 12466 19472 12478 19506
rect 13254 19472 13266 19506
rect 12466 19466 12830 19472
rect 12930 19466 13266 19472
rect 12388 19444 12434 19456
rect 12830 19453 12930 19463
rect 13298 19454 13344 19456
rect 12388 19276 12394 19444
rect 12428 19402 12434 19444
rect 13295 19444 13347 19454
rect 12428 19381 13295 19402
rect 12428 19329 12829 19381
rect 12929 19344 13295 19381
rect 12929 19329 13304 19344
rect 12428 19314 13304 19329
rect 12428 19276 12434 19314
rect 12388 19186 12434 19276
rect 13298 19276 13304 19314
rect 13338 19334 13347 19344
rect 13338 19276 13344 19334
rect 12478 19256 12678 19266
rect 12466 19208 12478 19254
rect 12678 19248 13266 19254
rect 13254 19214 13266 19248
rect 12678 19208 13266 19214
rect 12478 19194 12678 19204
rect 12388 19018 12394 19186
rect 12428 19145 12434 19186
rect 13298 19186 13344 19276
rect 13298 19145 13304 19186
rect 12428 19129 13304 19145
rect 12428 19077 12832 19129
rect 12932 19077 13304 19129
rect 12428 19057 13304 19077
rect 12428 19018 12434 19057
rect 12388 19006 12434 19018
rect 13298 19018 13304 19057
rect 13338 19018 13344 19186
rect 12830 18999 12930 19009
rect 13298 19006 13344 19018
rect 12466 18990 12830 18996
rect 12930 18990 13266 18996
rect 12466 18956 12478 18990
rect 13254 18956 13266 18990
rect 12466 18950 12830 18956
rect 12930 18950 13266 18956
rect 13521 18976 13573 19650
rect 12388 18928 12434 18940
rect 12830 18937 12930 18947
rect 13298 18938 13344 18940
rect 12388 18760 12394 18928
rect 12428 18893 12434 18928
rect 13295 18928 13347 18938
rect 12428 18805 13295 18893
rect 12428 18760 12434 18805
rect 13295 18788 13304 18802
rect 12388 18670 12434 18760
rect 13298 18760 13304 18788
rect 13338 18788 13347 18802
rect 13338 18760 13344 18788
rect 13054 18743 13254 18753
rect 12466 18732 13054 18738
rect 12466 18698 12478 18732
rect 12466 18692 13054 18698
rect 13254 18692 13266 18738
rect 13054 18677 13254 18687
rect 12388 18502 12394 18670
rect 12428 18634 12434 18670
rect 13298 18670 13344 18760
rect 13298 18634 13304 18670
rect 12428 18546 13304 18634
rect 12428 18502 12434 18546
rect 12388 18412 12434 18502
rect 13298 18502 13304 18546
rect 13338 18502 13344 18670
rect 12478 18489 12678 18499
rect 12466 18434 12478 18480
rect 12678 18474 13266 18480
rect 13254 18440 13266 18474
rect 12678 18434 13266 18440
rect 12478 18415 12678 18425
rect 12388 18244 12394 18412
rect 12428 18377 12434 18412
rect 13298 18412 13344 18502
rect 13298 18377 13304 18412
rect 12428 18289 13304 18377
rect 12428 18244 12434 18289
rect 12388 18154 12434 18244
rect 13298 18244 13304 18289
rect 13338 18244 13344 18412
rect 13054 18227 13254 18237
rect 12466 18216 13054 18222
rect 12466 18182 12478 18216
rect 12466 18176 13054 18182
rect 13254 18176 13266 18222
rect 13054 18161 13254 18171
rect 12388 17986 12394 18154
rect 12428 18121 12434 18154
rect 13298 18154 13344 18244
rect 13298 18121 13304 18154
rect 12428 18033 13304 18121
rect 12428 17986 12434 18033
rect 12388 17974 12434 17986
rect 13298 17986 13304 18033
rect 13338 17986 13344 18154
rect 12830 17967 12930 17977
rect 13298 17974 13344 17986
rect 13521 18202 13573 18876
rect 12466 17958 12830 17964
rect 12930 17958 13266 17964
rect 12466 17924 12478 17958
rect 13254 17924 13266 17958
rect 12466 17918 12830 17924
rect 12930 17918 13266 17924
rect 12388 17896 12434 17908
rect 12830 17905 12930 17915
rect 13298 17906 13344 17908
rect 12388 17728 12394 17896
rect 12428 17856 12434 17896
rect 13295 17896 13347 17906
rect 12428 17836 13295 17856
rect 12428 17784 12831 17836
rect 12931 17796 13295 17836
rect 12931 17784 13304 17796
rect 12428 17768 13304 17784
rect 12428 17728 12434 17768
rect 12388 17638 12434 17728
rect 13298 17728 13304 17768
rect 13338 17786 13347 17796
rect 13338 17728 13344 17786
rect 12478 17709 12678 17719
rect 12466 17660 12478 17706
rect 12678 17700 13266 17706
rect 13254 17666 13266 17700
rect 12678 17660 13266 17666
rect 12478 17647 12678 17657
rect 12388 17470 12394 17638
rect 12428 17599 12434 17638
rect 13298 17638 13344 17728
rect 13298 17599 13304 17638
rect 12428 17574 13304 17599
rect 12428 17522 12829 17574
rect 12929 17522 13304 17574
rect 12428 17506 13304 17522
rect 12428 17470 12434 17506
rect 12388 17458 12434 17470
rect 13298 17470 13304 17506
rect 13338 17470 13344 17638
rect 12830 17451 12930 17461
rect 13298 17458 13344 17470
rect 12466 17442 12830 17448
rect 12930 17442 13266 17448
rect 12466 17408 12478 17442
rect 13254 17408 13266 17442
rect 12466 17402 12830 17408
rect 12930 17402 13266 17408
rect 13521 17428 13573 18102
rect 12388 17380 12434 17392
rect 12830 17389 12930 17399
rect 13298 17390 13344 17392
rect 12388 17212 12394 17380
rect 12428 17341 12434 17380
rect 13295 17380 13347 17390
rect 12428 17254 13295 17341
rect 13347 17254 13357 17276
rect 12428 17253 13304 17254
rect 12428 17212 12434 17253
rect 13285 17231 13304 17253
rect 12388 17122 12434 17212
rect 13298 17212 13304 17231
rect 13338 17231 13357 17254
rect 13338 17212 13344 17231
rect 13054 17195 13254 17205
rect 12466 17184 13054 17190
rect 12466 17150 12478 17184
rect 12466 17144 13054 17150
rect 13254 17144 13266 17190
rect 13054 17129 13254 17139
rect 12388 16954 12394 17122
rect 12428 17082 12434 17122
rect 13298 17122 13344 17212
rect 13298 17082 13304 17122
rect 12428 16994 13304 17082
rect 12428 16954 12434 16994
rect 12388 16864 12434 16954
rect 13298 16954 13304 16994
rect 13338 16954 13344 17122
rect 12478 16941 12678 16951
rect 12466 16886 12478 16932
rect 12678 16926 13266 16932
rect 13254 16892 13266 16926
rect 12678 16886 13266 16892
rect 12478 16867 12678 16877
rect 12388 16696 12394 16864
rect 12428 16832 12434 16864
rect 13298 16864 13344 16954
rect 13298 16832 13304 16864
rect 12428 16744 13304 16832
rect 12428 16696 12434 16744
rect 12388 16606 12434 16696
rect 13298 16696 13304 16744
rect 13338 16696 13344 16864
rect 13054 16679 13254 16689
rect 12466 16668 13054 16674
rect 12466 16634 12478 16668
rect 12466 16628 13054 16634
rect 13254 16628 13266 16674
rect 13054 16613 13254 16623
rect 12388 16438 12394 16606
rect 12428 16569 12434 16606
rect 13298 16606 13344 16696
rect 13298 16569 13304 16606
rect 12428 16481 13304 16569
rect 12428 16438 12434 16481
rect 12388 16426 12434 16438
rect 13298 16438 13304 16481
rect 13338 16438 13344 16606
rect 12830 16419 12930 16429
rect 13298 16426 13344 16438
rect 13521 16654 13573 17328
rect 12466 16410 12830 16416
rect 12930 16410 13266 16416
rect 12466 16376 12478 16410
rect 13254 16376 13266 16410
rect 12466 16370 12830 16376
rect 12930 16370 13266 16376
rect 12388 16348 12434 16360
rect 12830 16357 12930 16367
rect 13298 16358 13344 16360
rect 12388 16180 12394 16348
rect 12428 16308 12434 16348
rect 13295 16348 13347 16358
rect 12428 16292 13295 16308
rect 12428 16240 12830 16292
rect 12930 16248 13295 16292
rect 12930 16240 13304 16248
rect 12428 16220 13304 16240
rect 12428 16180 12434 16220
rect 12388 16090 12434 16180
rect 13298 16180 13304 16220
rect 13338 16238 13347 16248
rect 13338 16180 13344 16238
rect 12478 16161 12678 16171
rect 12466 16112 12478 16158
rect 12678 16152 13266 16158
rect 13254 16118 13266 16152
rect 12678 16112 13266 16118
rect 12478 16099 12678 16109
rect 12388 15922 12394 16090
rect 12428 16045 12434 16090
rect 13298 16090 13344 16180
rect 13298 16045 13304 16090
rect 12428 16027 13304 16045
rect 12428 15975 12830 16027
rect 12930 15975 13304 16027
rect 12428 15956 13304 15975
rect 12428 15922 12434 15956
rect 12388 15910 12434 15922
rect 13298 15922 13304 15956
rect 13338 15922 13344 16090
rect 12830 15903 12930 15913
rect 13298 15910 13344 15922
rect 12466 15894 12830 15900
rect 12930 15894 13266 15900
rect 12466 15860 12478 15894
rect 13254 15860 13266 15894
rect 12466 15854 12830 15860
rect 12930 15854 13266 15860
rect 13521 15880 13573 16554
rect 12388 15832 12434 15844
rect 12830 15841 12930 15851
rect 13298 15842 13344 15844
rect 12388 15664 12394 15832
rect 12428 15796 12434 15832
rect 13295 15832 13347 15842
rect 12428 15732 13295 15796
rect 12428 15707 13304 15732
rect 12428 15664 12434 15707
rect 12388 15574 12434 15664
rect 13298 15664 13304 15707
rect 13338 15722 13347 15732
rect 13338 15664 13344 15722
rect 13054 15647 13254 15657
rect 12466 15636 13054 15642
rect 12466 15602 12478 15636
rect 12466 15596 13054 15602
rect 13254 15596 13266 15642
rect 13054 15581 13254 15591
rect 12388 15406 12394 15574
rect 12428 15532 12434 15574
rect 13298 15574 13344 15664
rect 13298 15532 13304 15574
rect 12428 15443 13304 15532
rect 12428 15406 12434 15443
rect 12388 15394 12434 15406
rect 13298 15406 13304 15443
rect 13338 15406 13344 15574
rect 12478 15393 12678 15403
rect 13298 15394 13344 15406
rect 12466 15338 12478 15384
rect 12678 15378 13266 15384
rect 13254 15344 13266 15378
rect 12678 15338 13266 15344
rect 12478 15319 12678 15329
rect 13521 15261 13573 15780
rect 13666 21556 13718 21566
rect 13947 21536 13959 21570
rect 13947 21530 14535 21536
rect 14735 21530 14747 21576
rect 13869 21518 13915 21520
rect 13666 21040 13718 21456
rect 13866 21508 13918 21518
rect 14535 21517 14735 21527
rect 14779 21508 14825 21520
rect 14779 21467 14785 21508
rect 13918 21447 14785 21467
rect 13918 21408 14258 21447
rect 13866 21398 13875 21408
rect 13869 21340 13875 21398
rect 13909 21395 14258 21408
rect 14358 21395 14785 21447
rect 13909 21379 14785 21395
rect 13909 21340 13915 21379
rect 13869 21328 13915 21340
rect 14779 21340 14785 21379
rect 14819 21340 14825 21508
rect 14260 21321 14360 21331
rect 14779 21328 14825 21340
rect 13947 21312 14260 21318
rect 14360 21312 14747 21318
rect 13947 21278 13959 21312
rect 14735 21278 14747 21312
rect 13947 21272 14260 21278
rect 14360 21272 14747 21278
rect 13869 21260 13915 21262
rect 13866 21250 13918 21260
rect 14260 21259 14360 21269
rect 14779 21250 14825 21262
rect 14779 21214 14785 21250
rect 13918 21126 14785 21214
rect 14779 21082 14785 21126
rect 14819 21082 14825 21250
rect 13866 21056 13918 21066
rect 14535 21065 14735 21075
rect 13666 20266 13718 20940
rect 13869 20992 13915 21056
rect 13947 21054 14535 21060
rect 13947 21020 13959 21054
rect 13947 21014 14535 21020
rect 14735 21014 14747 21060
rect 14535 20999 14735 21009
rect 13869 20824 13875 20992
rect 13909 20954 13915 20992
rect 14779 20992 14825 21082
rect 14779 20954 14785 20992
rect 13909 20866 14785 20954
rect 13909 20824 13915 20866
rect 13869 20734 13915 20824
rect 14779 20824 14785 20866
rect 14819 20824 14825 20992
rect 13959 20811 14159 20821
rect 13947 20756 13959 20802
rect 14159 20796 14747 20802
rect 14735 20762 14747 20796
rect 14159 20756 14747 20762
rect 13959 20737 14159 20747
rect 13869 20566 13875 20734
rect 13909 20695 13915 20734
rect 14779 20734 14825 20824
rect 14779 20695 14785 20734
rect 13909 20607 14785 20695
rect 13909 20566 13915 20607
rect 13869 20476 13915 20566
rect 14779 20566 14785 20607
rect 14819 20566 14825 20734
rect 14535 20549 14735 20559
rect 13947 20538 14535 20544
rect 13947 20504 13959 20538
rect 13947 20498 14535 20504
rect 14735 20498 14747 20544
rect 14535 20483 14735 20493
rect 13869 20308 13875 20476
rect 13909 20439 13915 20476
rect 14779 20476 14825 20566
rect 14779 20439 14785 20476
rect 13909 20351 14785 20439
rect 13909 20308 13915 20351
rect 13869 20296 13915 20308
rect 14779 20308 14785 20351
rect 14819 20308 14825 20476
rect 14260 20289 14360 20299
rect 14779 20296 14825 20308
rect 13947 20280 14260 20286
rect 14360 20280 14747 20286
rect 13947 20246 13959 20280
rect 14735 20246 14747 20280
rect 13947 20240 14260 20246
rect 14360 20240 14747 20246
rect 13869 20228 13915 20230
rect 13666 19492 13718 20166
rect 13866 20218 13918 20228
rect 14260 20227 14360 20237
rect 14779 20218 14825 20230
rect 14779 20187 14785 20218
rect 13918 20155 14785 20187
rect 13918 20118 14260 20155
rect 13866 20108 13875 20118
rect 13869 20050 13875 20108
rect 13909 20103 14260 20118
rect 14360 20103 14785 20155
rect 13909 20081 14785 20103
rect 13909 20050 13915 20081
rect 13869 19960 13915 20050
rect 14779 20050 14785 20081
rect 14819 20050 14825 20218
rect 14535 20031 14735 20041
rect 13947 20022 14535 20028
rect 13947 19988 13959 20022
rect 13947 19982 14535 19988
rect 14735 19982 14747 20028
rect 14535 19969 14735 19979
rect 13869 19792 13875 19960
rect 13909 19932 13915 19960
rect 14779 19960 14825 20050
rect 14779 19932 14785 19960
rect 13909 19900 14785 19932
rect 13909 19848 14262 19900
rect 14362 19848 14785 19900
rect 13909 19826 14785 19848
rect 13909 19792 13915 19826
rect 13869 19780 13915 19792
rect 14779 19792 14785 19826
rect 14819 19792 14825 19960
rect 14260 19773 14360 19783
rect 14779 19780 14825 19792
rect 13947 19764 14260 19770
rect 14360 19764 14747 19770
rect 13947 19730 13959 19764
rect 14735 19730 14747 19764
rect 13947 19724 14260 19730
rect 14360 19724 14747 19730
rect 13869 19712 13915 19714
rect 13866 19702 13918 19712
rect 14260 19711 14360 19721
rect 14779 19702 14825 19714
rect 14779 19659 14785 19702
rect 13918 19571 14785 19659
rect 14779 19534 14785 19571
rect 14819 19534 14825 19702
rect 13866 19508 13918 19518
rect 14535 19517 14735 19527
rect 13666 18718 13718 19392
rect 13869 19444 13915 19508
rect 13947 19506 14535 19512
rect 13947 19472 13959 19506
rect 13947 19466 14535 19472
rect 14735 19466 14747 19512
rect 14535 19451 14735 19461
rect 13869 19276 13875 19444
rect 13909 19404 13915 19444
rect 14779 19444 14825 19534
rect 14779 19404 14785 19444
rect 13909 19316 14785 19404
rect 13909 19276 13915 19316
rect 13869 19186 13915 19276
rect 14779 19276 14785 19316
rect 14819 19276 14825 19444
rect 13959 19263 14159 19273
rect 13947 19208 13959 19254
rect 14159 19248 14747 19254
rect 14735 19214 14747 19248
rect 14159 19208 14747 19214
rect 13959 19189 14159 19199
rect 13869 19018 13875 19186
rect 13909 19143 13915 19186
rect 14779 19186 14825 19276
rect 14779 19143 14785 19186
rect 13909 19055 14785 19143
rect 13909 19018 13915 19055
rect 13869 18928 13915 19018
rect 14779 19018 14785 19055
rect 14819 19018 14825 19186
rect 14535 19001 14735 19011
rect 13947 18990 14535 18996
rect 13947 18956 13959 18990
rect 13947 18950 14535 18956
rect 14735 18950 14747 18996
rect 14535 18935 14735 18945
rect 13869 18760 13875 18928
rect 13909 18887 13915 18928
rect 14779 18928 14825 19018
rect 14779 18887 14785 18928
rect 13909 18799 14785 18887
rect 13909 18760 13915 18799
rect 13869 18748 13915 18760
rect 14779 18760 14785 18799
rect 14819 18760 14825 18928
rect 14259 18741 14359 18751
rect 14779 18748 14825 18760
rect 13947 18732 14259 18738
rect 14359 18732 14747 18738
rect 13947 18698 13959 18732
rect 14735 18698 14747 18732
rect 13947 18692 14259 18698
rect 14359 18692 14747 18698
rect 13869 18680 13915 18682
rect 13666 17944 13718 18618
rect 13866 18670 13918 18680
rect 14259 18679 14359 18689
rect 14779 18670 14825 18682
rect 14779 18618 14785 18670
rect 13918 18604 14785 18618
rect 13918 18570 14262 18604
rect 13866 18560 13875 18570
rect 13869 18502 13875 18560
rect 13909 18552 14262 18570
rect 14362 18552 14785 18604
rect 13909 18537 14785 18552
rect 13909 18502 13915 18537
rect 13869 18412 13915 18502
rect 14779 18502 14785 18537
rect 14819 18502 14825 18670
rect 14535 18483 14735 18493
rect 13947 18474 14535 18480
rect 13947 18440 13959 18474
rect 13947 18434 14535 18440
rect 14735 18434 14747 18480
rect 14535 18421 14735 18431
rect 13869 18244 13875 18412
rect 13909 18358 13915 18412
rect 14779 18412 14825 18502
rect 14779 18358 14785 18412
rect 13909 18342 14785 18358
rect 13909 18290 14260 18342
rect 14360 18290 14785 18342
rect 13909 18277 14785 18290
rect 13909 18244 13915 18277
rect 13869 18232 13915 18244
rect 14779 18244 14785 18277
rect 14819 18244 14825 18412
rect 14260 18225 14360 18235
rect 14779 18232 14825 18244
rect 13947 18216 14260 18222
rect 14360 18216 14747 18222
rect 13947 18182 13959 18216
rect 14735 18182 14747 18216
rect 13947 18176 14260 18182
rect 14360 18176 14747 18182
rect 13869 18164 13915 18166
rect 13866 18154 13918 18164
rect 14260 18163 14360 18173
rect 14779 18154 14825 18166
rect 14779 18119 14785 18154
rect 13918 18031 14785 18119
rect 14779 17986 14785 18031
rect 14819 17986 14825 18154
rect 13866 17960 13918 17970
rect 14535 17969 14735 17979
rect 13666 17170 13718 17844
rect 13869 17896 13915 17960
rect 13947 17958 14535 17964
rect 13947 17924 13959 17958
rect 13947 17918 14535 17924
rect 14735 17918 14747 17964
rect 14535 17903 14735 17913
rect 13869 17728 13875 17896
rect 13909 17848 13915 17896
rect 14779 17896 14825 17986
rect 14779 17848 14785 17896
rect 13909 17760 14785 17848
rect 13909 17728 13915 17760
rect 13869 17638 13915 17728
rect 14779 17728 14785 17760
rect 14819 17728 14825 17896
rect 13959 17715 14159 17725
rect 13947 17660 13959 17706
rect 14159 17700 14747 17706
rect 14735 17666 14747 17700
rect 14159 17660 14747 17666
rect 13959 17641 14159 17651
rect 13869 17470 13875 17638
rect 13909 17596 13915 17638
rect 14779 17638 14825 17728
rect 14779 17596 14785 17638
rect 13909 17508 14785 17596
rect 13909 17470 13915 17508
rect 13869 17380 13915 17470
rect 14779 17470 14785 17508
rect 14819 17470 14825 17638
rect 14535 17453 14735 17463
rect 13947 17442 14535 17448
rect 13947 17408 13959 17442
rect 13947 17402 14535 17408
rect 14735 17402 14747 17448
rect 14535 17387 14735 17397
rect 13869 17212 13875 17380
rect 13909 17343 13915 17380
rect 14779 17380 14825 17470
rect 14779 17343 14785 17380
rect 13909 17255 14785 17343
rect 13909 17212 13915 17255
rect 13869 17200 13915 17212
rect 14779 17212 14785 17255
rect 14819 17212 14825 17380
rect 14260 17193 14360 17203
rect 14779 17200 14825 17212
rect 13947 17184 14260 17190
rect 14360 17184 14747 17190
rect 13947 17150 13959 17184
rect 14735 17150 14747 17184
rect 13947 17144 14260 17150
rect 14360 17144 14747 17150
rect 13869 17132 13915 17134
rect 13666 16396 13718 17070
rect 13866 17122 13918 17132
rect 14260 17131 14360 17141
rect 14779 17122 14825 17134
rect 14779 17076 14785 17122
rect 13918 17056 14785 17076
rect 13918 17022 14258 17056
rect 13866 17012 13875 17022
rect 13869 16954 13875 17012
rect 13909 17004 14258 17022
rect 14358 17004 14785 17056
rect 13909 16988 14785 17004
rect 13909 16954 13915 16988
rect 13869 16864 13915 16954
rect 14779 16954 14785 16988
rect 14819 16954 14825 17122
rect 14535 16935 14735 16945
rect 13947 16926 14535 16932
rect 13947 16892 13959 16926
rect 13947 16886 14535 16892
rect 14735 16886 14747 16932
rect 14535 16873 14735 16883
rect 13869 16696 13875 16864
rect 13909 16822 13915 16864
rect 14779 16864 14825 16954
rect 14779 16822 14785 16864
rect 13909 16800 14785 16822
rect 13909 16748 14259 16800
rect 14359 16748 14785 16800
rect 13909 16734 14785 16748
rect 13909 16696 13915 16734
rect 13869 16684 13915 16696
rect 14779 16696 14785 16734
rect 14819 16696 14825 16864
rect 14260 16677 14360 16687
rect 14779 16684 14825 16696
rect 13947 16668 14260 16674
rect 14360 16668 14747 16674
rect 13947 16634 13959 16668
rect 14735 16634 14747 16668
rect 13947 16628 14260 16634
rect 14360 16628 14747 16634
rect 13869 16616 13915 16618
rect 13866 16606 13918 16616
rect 14260 16615 14360 16625
rect 14779 16606 14825 16618
rect 14779 16559 14785 16606
rect 13918 16471 14785 16559
rect 14779 16438 14785 16471
rect 14819 16438 14825 16606
rect 14535 16421 14735 16431
rect 13866 16396 13918 16406
rect 13947 16410 14535 16416
rect 13666 15622 13718 16296
rect 13869 16348 13915 16396
rect 13947 16376 13959 16410
rect 13947 16370 14535 16376
rect 14735 16370 14747 16416
rect 14535 16355 14735 16365
rect 13869 16180 13875 16348
rect 13909 16310 13915 16348
rect 14779 16348 14825 16438
rect 14779 16310 14785 16348
rect 13909 16222 14785 16310
rect 13909 16180 13915 16222
rect 13869 16090 13915 16180
rect 14779 16180 14785 16222
rect 14819 16180 14825 16348
rect 13959 16167 14159 16177
rect 13947 16112 13959 16158
rect 14159 16152 14747 16158
rect 14735 16118 14747 16152
rect 14159 16112 14747 16118
rect 13959 16093 14159 16103
rect 13869 15922 13875 16090
rect 13909 16040 13915 16090
rect 14779 16090 14825 16180
rect 14779 16040 14785 16090
rect 13909 15952 14785 16040
rect 13909 15922 13915 15952
rect 13869 15832 13915 15922
rect 14779 15922 14785 15952
rect 14819 15922 14825 16090
rect 14534 15905 14734 15915
rect 13947 15894 14534 15900
rect 14734 15894 14747 15900
rect 13947 15860 13959 15894
rect 14735 15860 14747 15894
rect 13947 15854 14534 15860
rect 14734 15854 14747 15860
rect 14534 15839 14734 15849
rect 13869 15664 13875 15832
rect 13909 15791 13915 15832
rect 14779 15832 14825 15922
rect 14779 15791 14785 15832
rect 13909 15703 14785 15791
rect 13909 15664 13915 15703
rect 13869 15652 13915 15664
rect 14779 15664 14785 15703
rect 14819 15664 14825 15832
rect 14260 15645 14360 15655
rect 14779 15652 14825 15664
rect 13947 15636 14260 15642
rect 14360 15636 14747 15642
rect 13947 15602 13959 15636
rect 14735 15602 14747 15636
rect 13947 15596 14260 15602
rect 14360 15596 14747 15602
rect 13869 15584 13915 15586
rect 13666 15400 13718 15522
rect 13866 15574 13918 15584
rect 14260 15583 14360 15593
rect 14779 15574 14825 15586
rect 14779 15539 14785 15574
rect 13918 15522 14785 15539
rect 13918 15474 14262 15522
rect 13866 15464 13875 15474
rect 13869 15406 13875 15464
rect 13909 15470 14262 15474
rect 14362 15470 14785 15522
rect 13909 15451 14785 15470
rect 13909 15406 13915 15451
rect 13869 15394 13915 15406
rect 14779 15406 14785 15451
rect 14819 15406 14825 15574
rect 14535 15387 14735 15397
rect 14779 15394 14825 15406
rect 13947 15378 14535 15384
rect 13947 15344 13959 15378
rect 13947 15338 14535 15344
rect 14735 15338 14747 15384
rect 14535 15325 14735 15335
rect 14988 15315 14994 21656
rect 15106 15315 15112 21656
rect 15730 17060 15736 22467
rect 15927 17060 15933 22467
rect 16883 22449 17006 22459
rect 16871 22400 16883 22446
rect 17006 22440 17071 22446
rect 17059 22406 17071 22440
rect 17006 22400 17071 22406
rect 16096 22384 16156 22394
rect 16084 22335 16096 22381
rect 16212 22384 16272 22394
rect 16156 22375 16212 22381
rect 16156 22335 16212 22341
rect 16006 22313 16052 22325
rect 16096 22322 16156 22332
rect 16272 22335 16284 22381
rect 16784 22378 16830 22395
rect 16883 22387 17006 22397
rect 16212 22322 16272 22332
rect 16006 22145 16012 22313
rect 16046 22271 16052 22313
rect 16316 22313 16362 22325
rect 16316 22271 16322 22313
rect 16046 22204 16322 22271
rect 16046 22145 16052 22204
rect 16006 22123 16052 22145
rect 16316 22145 16322 22204
rect 16356 22145 16362 22313
rect 16316 22136 16362 22145
rect 16212 22126 16362 22136
rect 16006 22117 16212 22123
rect 16006 22083 16096 22117
rect 16006 22077 16212 22083
rect 16006 22055 16052 22077
rect 16272 22074 16362 22126
rect 16212 22064 16362 22074
rect 16006 21887 16012 22055
rect 16046 22004 16052 22055
rect 16316 22055 16362 22064
rect 16316 22004 16322 22055
rect 16046 21937 16322 22004
rect 16046 21887 16052 21937
rect 16006 21797 16052 21887
rect 16316 21887 16322 21937
rect 16356 21887 16362 22055
rect 16096 21868 16156 21878
rect 16084 21819 16096 21865
rect 16156 21859 16284 21865
rect 16272 21825 16284 21859
rect 16156 21819 16284 21825
rect 16096 21806 16156 21816
rect 16006 21629 16012 21797
rect 16046 21745 16052 21797
rect 16316 21797 16362 21887
rect 16316 21745 16322 21797
rect 16046 21678 16322 21745
rect 16046 21629 16052 21678
rect 16006 21607 16052 21629
rect 16316 21629 16322 21678
rect 16356 21629 16362 21797
rect 16316 21620 16362 21629
rect 16212 21610 16362 21620
rect 16006 21601 16212 21607
rect 16006 21567 16096 21601
rect 16006 21561 16212 21567
rect 16006 21539 16052 21561
rect 16272 21558 16362 21610
rect 16212 21548 16362 21558
rect 16006 21371 16012 21539
rect 16046 21485 16052 21539
rect 16316 21539 16362 21548
rect 16316 21485 16322 21539
rect 16046 21418 16322 21485
rect 16046 21371 16052 21418
rect 16006 21281 16052 21371
rect 16316 21371 16322 21418
rect 16356 21371 16362 21539
rect 16096 21352 16156 21362
rect 16084 21303 16096 21349
rect 16156 21343 16284 21349
rect 16272 21309 16284 21343
rect 16156 21303 16284 21309
rect 16096 21290 16156 21300
rect 16006 21113 16012 21281
rect 16046 21223 16052 21281
rect 16316 21281 16362 21371
rect 16316 21223 16322 21281
rect 16046 21156 16322 21223
rect 16046 21113 16052 21156
rect 16006 21101 16052 21113
rect 16316 21113 16322 21156
rect 16356 21113 16362 21281
rect 16096 21094 16156 21104
rect 16316 21101 16362 21113
rect 16784 22010 16790 22378
rect 16824 22341 16830 22378
rect 17112 22378 17158 22390
rect 17112 22341 17118 22378
rect 16824 22062 17118 22341
rect 16824 22010 16830 22062
rect 16784 21797 16830 22010
rect 17112 22010 17118 22062
rect 17152 22010 17158 22378
rect 16936 21991 17059 22001
rect 17112 21998 17158 22010
rect 16871 21982 16936 21988
rect 16871 21948 16883 21982
rect 16871 21942 16936 21948
rect 17059 21942 17071 21988
rect 16936 21929 17059 21939
rect 16883 21868 17006 21878
rect 16871 21819 16883 21865
rect 17006 21859 17071 21865
rect 17059 21825 17071 21859
rect 17006 21819 17071 21825
rect 16883 21806 17006 21816
rect 16784 21429 16790 21797
rect 16824 21765 16830 21797
rect 17112 21797 17158 21809
rect 17112 21765 17118 21797
rect 16824 21486 17118 21765
rect 16824 21429 16830 21486
rect 16084 21045 16096 21091
rect 16156 21085 16284 21091
rect 16272 21051 16284 21085
rect 16156 21045 16284 21051
rect 16006 21023 16052 21035
rect 16096 21032 16156 21042
rect 16006 20855 16012 21023
rect 16046 20963 16052 21023
rect 16316 21023 16362 21035
rect 16316 20963 16322 21023
rect 16046 20896 16322 20963
rect 16046 20855 16052 20896
rect 16006 20833 16052 20855
rect 16316 20855 16322 20896
rect 16356 20855 16362 21023
rect 16316 20846 16362 20855
rect 16212 20836 16362 20846
rect 16006 20827 16212 20833
rect 16006 20793 16096 20827
rect 16006 20787 16212 20793
rect 16006 20765 16052 20787
rect 16272 20784 16362 20836
rect 16212 20774 16362 20784
rect 16006 20597 16012 20765
rect 16046 20713 16052 20765
rect 16316 20765 16362 20774
rect 16316 20713 16322 20765
rect 16046 20646 16322 20713
rect 16046 20597 16052 20646
rect 16006 20507 16052 20597
rect 16316 20597 16322 20646
rect 16356 20597 16362 20765
rect 16096 20578 16156 20588
rect 16084 20529 16096 20575
rect 16156 20569 16284 20575
rect 16272 20535 16284 20569
rect 16156 20529 16284 20535
rect 16096 20516 16156 20526
rect 16006 20339 16012 20507
rect 16046 20454 16052 20507
rect 16316 20507 16362 20597
rect 16316 20454 16322 20507
rect 16046 20387 16322 20454
rect 16046 20339 16052 20387
rect 16006 20317 16052 20339
rect 16316 20339 16322 20387
rect 16356 20339 16362 20507
rect 16316 20330 16362 20339
rect 16212 20320 16362 20330
rect 16006 20311 16212 20317
rect 16006 20277 16096 20311
rect 16006 20271 16212 20277
rect 16006 20249 16052 20271
rect 16272 20268 16362 20320
rect 16212 20258 16362 20268
rect 16006 20081 16012 20249
rect 16046 20193 16052 20249
rect 16316 20249 16362 20258
rect 16316 20193 16322 20249
rect 16046 20126 16322 20193
rect 16046 20081 16052 20126
rect 16006 19991 16052 20081
rect 16316 20081 16322 20126
rect 16356 20081 16362 20249
rect 16096 20062 16156 20072
rect 16084 20013 16096 20059
rect 16156 20053 16284 20059
rect 16272 20019 16284 20053
rect 16156 20013 16284 20019
rect 16096 20000 16156 20010
rect 16006 19823 16012 19991
rect 16046 19936 16052 19991
rect 16316 19991 16362 20081
rect 16316 19936 16322 19991
rect 16046 19869 16322 19936
rect 16046 19823 16052 19869
rect 16006 19811 16052 19823
rect 16316 19823 16322 19869
rect 16356 19823 16362 19991
rect 16096 19804 16156 19814
rect 16316 19811 16362 19823
rect 16784 20507 16830 21429
rect 17112 21429 17118 21486
rect 17152 21429 17158 21797
rect 16935 21410 17059 21420
rect 17112 21417 17158 21429
rect 16871 21401 16935 21407
rect 16871 21367 16883 21401
rect 16871 21361 16935 21367
rect 17059 21361 17071 21407
rect 16935 21348 17059 21358
rect 17320 21170 17324 21228
rect 16883 20578 16996 20588
rect 16871 20529 16883 20575
rect 16996 20569 17071 20575
rect 17059 20535 17071 20569
rect 16996 20529 17071 20535
rect 16883 20516 16996 20526
rect 16784 20139 16790 20507
rect 16824 20455 16830 20507
rect 17112 20507 17158 20519
rect 17112 20455 17118 20507
rect 16824 20176 17118 20455
rect 16824 20139 16830 20176
rect 16084 19755 16096 19801
rect 16156 19795 16284 19801
rect 16272 19761 16284 19795
rect 16156 19755 16284 19761
rect 16006 19733 16052 19745
rect 16096 19742 16156 19752
rect 16006 19565 16012 19733
rect 16046 19678 16052 19733
rect 16316 19733 16362 19745
rect 16316 19678 16322 19733
rect 16046 19611 16322 19678
rect 16046 19565 16052 19611
rect 16006 19543 16052 19565
rect 16316 19565 16322 19611
rect 16356 19565 16362 19733
rect 16316 19556 16362 19565
rect 16212 19546 16362 19556
rect 16006 19537 16212 19543
rect 16006 19503 16096 19537
rect 16006 19497 16212 19503
rect 16006 19475 16052 19497
rect 16272 19494 16362 19546
rect 16212 19484 16362 19494
rect 16006 19307 16012 19475
rect 16046 19416 16052 19475
rect 16316 19475 16362 19484
rect 16316 19416 16322 19475
rect 16046 19349 16322 19416
rect 16046 19307 16052 19349
rect 16006 19217 16052 19307
rect 16316 19307 16322 19349
rect 16356 19307 16362 19475
rect 16096 19288 16156 19298
rect 16084 19239 16096 19285
rect 16156 19279 16284 19285
rect 16272 19245 16284 19279
rect 16156 19239 16284 19245
rect 16096 19226 16156 19236
rect 16006 19049 16012 19217
rect 16046 19163 16052 19217
rect 16316 19217 16362 19307
rect 16316 19163 16322 19217
rect 16046 19096 16322 19163
rect 16046 19049 16052 19096
rect 16006 19027 16052 19049
rect 16316 19049 16322 19096
rect 16356 19049 16362 19217
rect 16316 19040 16362 19049
rect 16212 19030 16362 19040
rect 16006 19021 16212 19027
rect 16006 18987 16096 19021
rect 16006 18981 16212 18987
rect 16006 18959 16052 18981
rect 16272 18978 16362 19030
rect 16212 18968 16362 18978
rect 16006 18791 16012 18959
rect 16046 18902 16052 18959
rect 16316 18959 16362 18968
rect 16316 18902 16322 18959
rect 16046 18835 16322 18902
rect 16046 18791 16052 18835
rect 16006 18701 16052 18791
rect 16316 18791 16322 18835
rect 16356 18791 16362 18959
rect 16096 18772 16156 18782
rect 16084 18723 16096 18769
rect 16156 18763 16284 18769
rect 16272 18729 16284 18763
rect 16156 18723 16284 18729
rect 16096 18710 16156 18720
rect 16006 18533 16012 18701
rect 16046 18648 16052 18701
rect 16316 18701 16362 18791
rect 16316 18648 16322 18701
rect 16046 18581 16322 18648
rect 16046 18533 16052 18581
rect 16006 18521 16052 18533
rect 16316 18533 16322 18581
rect 16356 18533 16362 18701
rect 16096 18514 16156 18524
rect 16316 18521 16362 18533
rect 16784 19217 16830 20139
rect 17112 20139 17118 20176
rect 17152 20139 17158 20507
rect 16936 20120 17059 20130
rect 17112 20127 17158 20139
rect 16871 20111 16936 20117
rect 16871 20077 16883 20111
rect 16871 20071 16936 20077
rect 17059 20071 17071 20117
rect 16936 20058 17059 20068
rect 16883 19288 16996 19298
rect 16871 19239 16883 19285
rect 16996 19279 17071 19285
rect 17059 19245 17071 19279
rect 16996 19239 17071 19245
rect 16883 19226 16996 19236
rect 16784 18849 16790 19217
rect 16824 19174 16830 19217
rect 17112 19217 17158 19229
rect 17112 19174 17118 19217
rect 16824 18895 17118 19174
rect 16824 18849 16830 18895
rect 16084 18465 16096 18511
rect 16156 18505 16284 18511
rect 16272 18471 16284 18505
rect 16156 18465 16284 18471
rect 16006 18443 16052 18455
rect 16096 18452 16156 18462
rect 16006 18275 16012 18443
rect 16046 18396 16052 18443
rect 16316 18443 16362 18455
rect 16316 18396 16322 18443
rect 16046 18329 16322 18396
rect 16046 18275 16052 18329
rect 16006 18253 16052 18275
rect 16316 18275 16322 18329
rect 16356 18275 16362 18443
rect 16316 18266 16362 18275
rect 16212 18256 16362 18266
rect 16006 18247 16212 18253
rect 16006 18213 16096 18247
rect 16006 18207 16212 18213
rect 16006 18185 16052 18207
rect 16272 18204 16362 18256
rect 16212 18194 16362 18204
rect 16006 18017 16012 18185
rect 16046 18136 16052 18185
rect 16316 18185 16362 18194
rect 16316 18136 16322 18185
rect 16046 18069 16322 18136
rect 16046 18017 16052 18069
rect 16006 17927 16052 18017
rect 16316 18017 16322 18069
rect 16356 18017 16362 18185
rect 16096 17998 16156 18008
rect 16084 17949 16096 17995
rect 16156 17989 16284 17995
rect 16272 17955 16284 17989
rect 16156 17949 16284 17955
rect 16096 17936 16156 17946
rect 16006 17759 16012 17927
rect 16046 17879 16052 17927
rect 16316 17927 16362 18017
rect 16316 17879 16322 17927
rect 16046 17812 16322 17879
rect 16046 17759 16052 17812
rect 16006 17737 16052 17759
rect 16316 17759 16322 17812
rect 16356 17759 16362 17927
rect 16316 17750 16362 17759
rect 16212 17740 16362 17750
rect 16006 17731 16212 17737
rect 16006 17697 16096 17731
rect 16006 17691 16212 17697
rect 16006 17669 16052 17691
rect 16272 17688 16362 17740
rect 16212 17678 16362 17688
rect 16006 17501 16012 17669
rect 16046 17617 16052 17669
rect 16316 17669 16362 17678
rect 16316 17617 16322 17669
rect 16046 17550 16322 17617
rect 16046 17501 16052 17550
rect 16006 17411 16052 17501
rect 16316 17501 16322 17550
rect 16356 17501 16362 17669
rect 16096 17482 16156 17492
rect 16084 17433 16096 17479
rect 16156 17473 16284 17479
rect 16272 17439 16284 17473
rect 16156 17433 16284 17439
rect 16096 17420 16156 17430
rect 16006 17243 16012 17411
rect 16046 17359 16052 17411
rect 16316 17411 16362 17501
rect 16316 17359 16322 17411
rect 16046 17292 16322 17359
rect 16046 17243 16052 17292
rect 16006 17231 16052 17243
rect 16316 17243 16322 17292
rect 16356 17243 16362 17411
rect 16096 17224 16156 17234
rect 16316 17231 16362 17243
rect 16784 17927 16830 18849
rect 17112 18849 17118 18895
rect 17152 18849 17158 19217
rect 16936 18830 17059 18840
rect 17112 18837 17158 18849
rect 16871 18821 16936 18827
rect 16871 18787 16883 18821
rect 16871 18781 16936 18787
rect 17059 18781 17071 18827
rect 16936 18768 17059 18778
rect 16883 17998 16996 18008
rect 16871 17949 16883 17995
rect 16996 17989 17071 17995
rect 17059 17955 17071 17989
rect 16996 17949 17071 17955
rect 16883 17936 16996 17946
rect 16784 17559 16790 17927
rect 16824 17876 16830 17927
rect 17112 17927 17158 17939
rect 17112 17876 17118 17927
rect 16824 17597 17118 17876
rect 16824 17559 16830 17597
rect 16084 17175 16096 17221
rect 16156 17215 16284 17221
rect 16272 17181 16284 17215
rect 16156 17175 16284 17181
rect 16096 17162 16156 17172
rect 15730 17048 15933 17060
rect 16784 16839 16830 17559
rect 17112 17559 17118 17597
rect 17152 17559 17158 17927
rect 16936 17540 17059 17550
rect 17112 17547 17158 17559
rect 16871 17531 16936 17537
rect 16871 17497 16883 17531
rect 16871 17491 16936 17497
rect 17059 17491 17071 17537
rect 16936 17478 17059 17488
rect 17324 17490 17330 21143
rect 22056 21625 22066 23052
rect 23409 22876 23955 22882
rect 23409 22875 23419 22876
rect 22404 21872 22414 22875
rect 23323 22756 23333 22766
rect 22654 22750 23333 22756
rect 23742 22756 23752 22766
rect 22654 22716 22666 22750
rect 22654 22710 23333 22716
rect 23323 22701 23333 22710
rect 23742 22710 23754 22756
rect 23742 22701 23752 22710
rect 22576 22688 22622 22700
rect 22576 22673 22582 22688
rect 22616 22673 22622 22688
rect 23786 22688 23832 22700
rect 22561 22533 22571 22673
rect 22627 22621 22637 22673
rect 23786 22621 23792 22688
rect 22627 22533 23792 22621
rect 22576 22420 22582 22533
rect 22616 22460 23792 22533
rect 22616 22420 22622 22460
rect 22576 22330 22622 22420
rect 23786 22420 23792 22460
rect 23826 22420 23832 22688
rect 22656 22398 22666 22407
rect 22654 22352 22666 22398
rect 23166 22398 23176 22407
rect 23166 22392 23754 22398
rect 23742 22358 23754 22392
rect 22656 22343 22666 22352
rect 23166 22352 23754 22358
rect 23166 22343 23176 22352
rect 22576 22062 22582 22330
rect 22616 22266 22622 22330
rect 23786 22330 23832 22420
rect 23786 22266 23792 22330
rect 22616 22105 23792 22266
rect 22616 22062 22622 22105
rect 22576 22050 22622 22062
rect 23786 22062 23792 22105
rect 23826 22062 23832 22330
rect 23786 22050 23832 22062
rect 23323 22040 23333 22050
rect 22654 22034 23333 22040
rect 23742 22040 23752 22050
rect 22654 22000 22666 22034
rect 22654 21994 23333 22000
rect 23323 21985 23333 21994
rect 23742 21994 23754 22040
rect 23742 21985 23752 21994
rect 23945 21872 23955 22876
rect 22404 21866 23955 21872
rect 24731 22882 24737 23222
rect 24897 23006 24907 23008
rect 24895 22956 24907 23006
rect 25109 23006 25119 23008
rect 25731 23006 25741 23007
rect 25109 23000 25316 23006
rect 25304 22962 25316 23000
rect 25109 22956 25316 22962
rect 25534 23000 25741 23006
rect 25943 23006 25953 23007
rect 25534 22962 25546 23000
rect 25534 22956 25741 22962
rect 25731 22955 25741 22956
rect 25943 22956 25955 23006
rect 25943 22955 25953 22956
rect 24166 22876 24737 22882
rect 22293 21625 23955 21627
rect 22060 21621 23955 21625
rect 22060 21613 22299 21621
rect 23945 21616 23955 21621
rect 24166 21616 24176 22876
rect 24536 22870 24737 22876
rect 23949 21604 24172 21616
rect 17475 21170 17479 21228
rect 17469 17490 17475 21143
rect 17324 17478 17475 17490
rect 17210 17028 17357 17040
rect 16883 16916 17023 16926
rect 16871 16861 16883 16907
rect 17023 16901 17071 16907
rect 17059 16867 17071 16901
rect 17023 16861 17071 16867
rect 16883 16842 17023 16852
rect 16784 16671 16790 16839
rect 16824 16814 16830 16839
rect 17112 16839 17158 16851
rect 17112 16814 17118 16839
rect 16824 16696 17118 16814
rect 16824 16671 16830 16696
rect 16784 16581 16830 16671
rect 17112 16671 17118 16696
rect 17152 16671 17158 16839
rect 16919 16652 17059 16662
rect 17112 16659 17158 16671
rect 16871 16643 16919 16649
rect 16871 16609 16883 16643
rect 16871 16603 16919 16609
rect 17059 16603 17071 16649
rect 16919 16590 17059 16600
rect 16784 16413 16790 16581
rect 16824 16562 16830 16581
rect 17112 16581 17158 16593
rect 17112 16562 17118 16581
rect 16824 16444 17118 16562
rect 16824 16413 16830 16444
rect 15334 16322 16377 16326
rect 15322 16316 16389 16322
rect 15322 16208 15334 16316
rect 16377 16208 16389 16316
rect 15322 16202 16389 16208
rect 15334 16198 16377 16202
rect 16784 16182 16830 16413
rect 17112 16413 17118 16444
rect 17152 16413 17158 16581
rect 16883 16400 17023 16410
rect 17112 16401 17158 16413
rect 16871 16345 16883 16391
rect 17023 16385 17071 16391
rect 17059 16351 17071 16385
rect 17023 16345 17071 16351
rect 16883 16326 17023 16336
rect 16784 16176 16971 16182
rect 16784 16142 16883 16176
rect 16959 16142 16971 16176
rect 16784 16136 16971 16142
rect 16784 16118 16830 16136
rect 16763 16114 16830 16118
rect 16763 16108 16790 16114
rect 16824 16108 16830 16114
rect 16338 16083 16498 16095
rect 15575 16015 16185 16053
rect 15575 15941 15580 16015
rect 16180 15941 16185 16015
rect 15575 15908 16185 15941
rect 15575 15874 15620 15908
rect 15654 15874 15720 15908
rect 15754 15874 15820 15908
rect 15854 15874 15920 15908
rect 15954 15874 16020 15908
rect 16054 15874 16120 15908
rect 16154 15874 16185 15908
rect 14988 15302 15112 15315
rect 15149 15834 15257 15846
rect 15149 15307 15155 15834
rect 15251 15307 15257 15834
rect 15149 15295 15257 15307
rect 15575 15808 16185 15874
rect 15575 15774 15620 15808
rect 15654 15774 15720 15808
rect 15754 15774 15820 15808
rect 15854 15774 15920 15808
rect 15954 15774 16020 15808
rect 16054 15774 16120 15808
rect 16154 15774 16185 15808
rect 15575 15708 16185 15774
rect 15575 15674 15620 15708
rect 15654 15674 15720 15708
rect 15754 15674 15820 15708
rect 15854 15674 15920 15708
rect 15954 15674 16020 15708
rect 16054 15674 16120 15708
rect 16154 15674 16185 15708
rect 15575 15608 16185 15674
rect 15575 15574 15620 15608
rect 15654 15574 15720 15608
rect 15754 15574 15820 15608
rect 15854 15574 15920 15608
rect 15954 15574 16020 15608
rect 16054 15574 16120 15608
rect 16154 15574 16185 15608
rect 15575 15508 16185 15574
rect 15575 15474 15620 15508
rect 15654 15474 15720 15508
rect 15754 15474 15820 15508
rect 15854 15474 15920 15508
rect 15954 15474 16020 15508
rect 16054 15474 16120 15508
rect 16154 15474 16185 15508
rect 15575 15443 16185 15474
rect 15575 15261 15627 15443
rect 15767 15287 16246 15291
rect 13521 15209 15627 15261
rect 15755 15281 16258 15287
rect 12309 15185 12461 15189
rect 13299 15185 13447 15189
rect 12047 15110 12233 15122
rect 12297 15179 12473 15185
rect 12297 15125 12309 15179
rect 12461 15125 12473 15179
rect 12297 15119 12473 15125
rect 13287 15179 13459 15185
rect 13287 15125 13299 15179
rect 13447 15125 13459 15179
rect 15755 15161 15767 15281
rect 16246 15161 16258 15281
rect 16338 15258 16344 16083
rect 16492 15258 16498 16083
rect 16828 16064 16830 16108
rect 17012 16114 17058 16126
rect 17012 16064 17018 16114
rect 16828 15782 17018 16064
rect 16828 15749 16830 15782
rect 16763 15746 16790 15749
rect 16824 15746 16830 15749
rect 16763 15739 16830 15746
rect 16784 15664 16830 15739
rect 17012 15746 17018 15782
rect 17052 15746 17058 16114
rect 17210 16042 17216 17028
rect 17351 16042 17357 17028
rect 17210 16030 17218 16042
rect 16883 15727 16959 15737
rect 17012 15734 17058 15746
rect 16871 15678 16883 15724
rect 16959 15678 16971 15724
rect 16883 15665 16959 15675
rect 16763 15656 16830 15664
rect 16763 15654 16790 15656
rect 16824 15654 16830 15656
rect 16828 15617 16830 15654
rect 17012 15656 17058 15668
rect 17012 15617 17018 15656
rect 16828 15335 17018 15617
rect 16828 15295 16830 15335
rect 16763 15288 16790 15295
rect 16824 15288 16830 15295
rect 16763 15285 16830 15288
rect 16338 15246 16498 15258
rect 16784 15266 16830 15285
rect 17012 15288 17018 15335
rect 17052 15288 17058 15656
rect 17012 15276 17058 15288
rect 16784 15260 16971 15266
rect 16784 15226 16883 15260
rect 16959 15226 16971 15260
rect 16784 15220 16971 15226
rect 15755 15155 16258 15161
rect 15767 15151 16246 15155
rect 13287 15119 13459 15125
rect 12309 15115 12461 15119
rect 13299 15115 13447 15119
rect 17212 15049 17218 16030
rect 17350 16030 17357 16042
rect 17423 17029 17583 17041
rect 17350 15049 17356 16030
rect 17212 15037 17356 15049
rect 17423 15050 17429 17029
rect 17577 15050 17583 17029
rect 17423 15038 17583 15050
rect 17898 11104 25720 11110
rect 17898 11015 17910 11104
rect 25708 11015 25720 11104
rect 17898 11009 25720 11015
rect 18028 10747 25475 10753
rect 18028 10713 18237 10747
rect 21805 10713 21895 10747
rect 25463 10713 25475 10747
rect 18028 10707 25475 10713
rect 18028 10654 18228 10707
rect 7847 10480 7991 10492
rect 2682 10407 2868 10419
rect 2944 10410 3096 10414
rect 3934 10410 4082 10414
rect 2682 3829 2688 10407
rect 2862 3829 2868 10407
rect 2932 10404 3108 10410
rect 2932 10350 2944 10404
rect 3096 10350 3108 10404
rect 2932 10344 3108 10350
rect 3922 10404 4094 10410
rect 3922 10350 3934 10404
rect 4082 10350 4094 10404
rect 6402 10374 6881 10378
rect 3922 10344 4094 10350
rect 6390 10368 6893 10374
rect 2944 10340 3096 10344
rect 3934 10340 4082 10344
rect 4156 10268 6262 10320
rect 3113 10200 3313 10210
rect 3101 10145 3113 10191
rect 3313 10185 3901 10191
rect 3889 10151 3901 10185
rect 3313 10145 3901 10151
rect 3023 10123 3069 10135
rect 3113 10126 3313 10136
rect 3023 9955 3029 10123
rect 3063 10086 3069 10123
rect 3933 10123 3979 10135
rect 3933 10086 3939 10123
rect 3063 9997 3939 10086
rect 3063 9955 3069 9997
rect 3023 9865 3069 9955
rect 3933 9955 3939 9997
rect 3973 9955 3979 10123
rect 3689 9938 3889 9948
rect 3101 9927 3689 9933
rect 3101 9893 3113 9927
rect 3101 9887 3689 9893
rect 3889 9887 3901 9933
rect 3689 9872 3889 9882
rect 3023 9697 3029 9865
rect 3063 9822 3069 9865
rect 3933 9865 3979 9955
rect 3933 9822 3939 9865
rect 3063 9797 3939 9822
rect 3973 9807 3979 9865
rect 3973 9797 3982 9807
rect 3063 9733 3930 9797
rect 3063 9697 3069 9733
rect 3023 9685 3069 9697
rect 3465 9678 3565 9688
rect 3930 9687 3982 9697
rect 4156 9749 4208 10268
rect 5623 10214 5747 10227
rect 5170 10194 5370 10204
rect 4582 10185 5170 10191
rect 4582 10151 4594 10185
rect 4582 10145 5170 10151
rect 5370 10145 5382 10191
rect 3933 9685 3979 9687
rect 3101 9669 3465 9675
rect 3565 9669 3901 9675
rect 3101 9635 3113 9669
rect 3889 9635 3901 9669
rect 3101 9629 3465 9635
rect 3565 9629 3901 9635
rect 3023 9607 3069 9619
rect 3465 9616 3565 9626
rect 3023 9439 3029 9607
rect 3063 9573 3069 9607
rect 3933 9607 3979 9619
rect 3933 9573 3939 9607
rect 3063 9554 3939 9573
rect 3063 9502 3465 9554
rect 3565 9502 3939 9554
rect 3063 9484 3939 9502
rect 3063 9439 3069 9484
rect 3023 9349 3069 9439
rect 3933 9439 3939 9484
rect 3973 9439 3979 9607
rect 3113 9420 3313 9430
rect 3101 9371 3113 9417
rect 3313 9411 3901 9417
rect 3889 9377 3901 9411
rect 3313 9371 3901 9377
rect 3113 9358 3313 9368
rect 3023 9181 3029 9349
rect 3063 9309 3069 9349
rect 3933 9349 3979 9439
rect 3933 9309 3939 9349
rect 3063 9289 3939 9309
rect 3063 9237 3465 9289
rect 3565 9281 3939 9289
rect 3973 9291 3979 9349
rect 3973 9281 3982 9291
rect 3565 9237 3930 9281
rect 3063 9221 3930 9237
rect 3063 9181 3069 9221
rect 3023 9169 3069 9181
rect 3465 9162 3565 9172
rect 3930 9171 3982 9181
rect 3933 9169 3979 9171
rect 3101 9153 3465 9159
rect 3565 9153 3901 9159
rect 3101 9119 3113 9153
rect 3889 9119 3901 9153
rect 3101 9113 3465 9119
rect 3565 9113 3901 9119
rect 3023 9091 3069 9103
rect 3465 9100 3565 9110
rect 3023 8923 3029 9091
rect 3063 9048 3069 9091
rect 3933 9091 3979 9103
rect 3933 9048 3939 9091
rect 3063 8960 3939 9048
rect 3063 8923 3069 8960
rect 3023 8833 3069 8923
rect 3933 8923 3939 8960
rect 3973 8923 3979 9091
rect 3689 8906 3889 8916
rect 3101 8895 3689 8901
rect 3101 8861 3113 8895
rect 3101 8855 3689 8861
rect 3889 8855 3901 8901
rect 3689 8840 3889 8850
rect 3023 8665 3029 8833
rect 3063 8785 3069 8833
rect 3933 8833 3979 8923
rect 3933 8785 3939 8833
rect 3063 8697 3939 8785
rect 3063 8665 3069 8697
rect 3023 8575 3069 8665
rect 3933 8665 3939 8697
rect 3973 8665 3979 8833
rect 3113 8652 3313 8662
rect 3101 8597 3113 8643
rect 3313 8637 3901 8643
rect 3889 8603 3901 8637
rect 3313 8597 3901 8603
rect 3113 8578 3313 8588
rect 3023 8407 3029 8575
rect 3063 8535 3069 8575
rect 3933 8575 3979 8665
rect 3933 8535 3939 8575
rect 3063 8447 3939 8535
rect 3063 8407 3069 8447
rect 3023 8317 3069 8407
rect 3933 8407 3939 8447
rect 3973 8407 3979 8575
rect 3689 8390 3889 8400
rect 3101 8379 3689 8385
rect 3101 8345 3113 8379
rect 3101 8339 3689 8345
rect 3889 8339 3901 8385
rect 3689 8324 3889 8334
rect 3023 8149 3029 8317
rect 3063 8276 3069 8317
rect 3933 8317 3979 8407
rect 3933 8298 3939 8317
rect 3920 8276 3939 8298
rect 3063 8275 3939 8276
rect 3973 8298 3979 8317
rect 4156 8975 4208 9649
rect 3973 8275 3992 8298
rect 3063 8188 3930 8275
rect 3063 8149 3069 8188
rect 3023 8137 3069 8149
rect 3982 8253 3992 8275
rect 3465 8130 3565 8140
rect 3930 8139 3982 8149
rect 4156 8201 4208 8875
rect 3933 8137 3979 8139
rect 3101 8121 3465 8127
rect 3565 8121 3901 8127
rect 3101 8087 3113 8121
rect 3889 8087 3901 8121
rect 3101 8081 3465 8087
rect 3565 8081 3901 8087
rect 3023 8059 3069 8071
rect 3465 8068 3565 8078
rect 3023 7891 3029 8059
rect 3063 8023 3069 8059
rect 3933 8059 3979 8071
rect 3933 8023 3939 8059
rect 3063 8007 3939 8023
rect 3063 7955 3464 8007
rect 3564 7955 3939 8007
rect 3063 7930 3939 7955
rect 3063 7891 3069 7930
rect 3023 7801 3069 7891
rect 3933 7891 3939 7930
rect 3973 7891 3979 8059
rect 3113 7872 3313 7882
rect 3101 7823 3113 7869
rect 3313 7863 3901 7869
rect 3889 7829 3901 7863
rect 3313 7823 3901 7829
rect 3113 7810 3313 7820
rect 3023 7633 3029 7801
rect 3063 7761 3069 7801
rect 3933 7801 3979 7891
rect 3933 7761 3939 7801
rect 3063 7745 3939 7761
rect 3063 7693 3466 7745
rect 3566 7733 3939 7745
rect 3973 7743 3979 7801
rect 3973 7733 3982 7743
rect 3566 7693 3930 7733
rect 3063 7673 3930 7693
rect 3063 7633 3069 7673
rect 3023 7621 3069 7633
rect 3465 7614 3565 7624
rect 3930 7623 3982 7633
rect 3933 7621 3979 7623
rect 3101 7605 3465 7611
rect 3565 7605 3901 7611
rect 3101 7571 3113 7605
rect 3889 7571 3901 7605
rect 3101 7565 3465 7571
rect 3565 7565 3901 7571
rect 3023 7543 3069 7555
rect 3465 7552 3565 7562
rect 3023 7375 3029 7543
rect 3063 7496 3069 7543
rect 3933 7543 3979 7555
rect 3933 7496 3939 7543
rect 3063 7408 3939 7496
rect 3063 7375 3069 7408
rect 3023 7285 3069 7375
rect 3933 7375 3939 7408
rect 3973 7375 3979 7543
rect 3689 7358 3889 7368
rect 3101 7347 3689 7353
rect 3101 7313 3113 7347
rect 3101 7307 3689 7313
rect 3889 7307 3901 7353
rect 3689 7292 3889 7302
rect 3023 7117 3029 7285
rect 3063 7240 3069 7285
rect 3933 7285 3979 7375
rect 3933 7240 3939 7285
rect 3063 7152 3939 7240
rect 3063 7117 3069 7152
rect 3023 7027 3069 7117
rect 3933 7117 3939 7152
rect 3973 7117 3979 7285
rect 3113 7104 3313 7114
rect 3101 7049 3113 7095
rect 3313 7089 3901 7095
rect 3889 7055 3901 7089
rect 3313 7049 3901 7055
rect 3113 7030 3313 7040
rect 3023 6859 3029 7027
rect 3063 6983 3069 7027
rect 3933 7027 3979 7117
rect 3933 6983 3939 7027
rect 3063 6895 3939 6983
rect 3063 6859 3069 6895
rect 3023 6769 3069 6859
rect 3933 6859 3939 6895
rect 3973 6859 3979 7027
rect 3689 6842 3889 6852
rect 3101 6831 3689 6837
rect 3101 6797 3113 6831
rect 3101 6791 3689 6797
rect 3889 6791 3901 6837
rect 3689 6776 3889 6786
rect 3023 6601 3029 6769
rect 3063 6724 3069 6769
rect 3933 6769 3979 6859
rect 3933 6741 3939 6769
rect 3930 6727 3939 6741
rect 3973 6741 3979 6769
rect 4156 7427 4208 8101
rect 3973 6727 3982 6741
rect 3063 6636 3930 6724
rect 3063 6601 3069 6636
rect 3023 6589 3069 6601
rect 3465 6582 3565 6592
rect 3930 6591 3982 6601
rect 4156 6653 4208 7327
rect 3933 6589 3979 6591
rect 3101 6573 3465 6579
rect 3565 6573 3901 6579
rect 3101 6539 3113 6573
rect 3889 6539 3901 6573
rect 3101 6533 3465 6539
rect 3565 6533 3901 6539
rect 3023 6511 3069 6523
rect 3465 6520 3565 6530
rect 3023 6343 3029 6511
rect 3063 6472 3069 6511
rect 3933 6511 3979 6523
rect 3933 6472 3939 6511
rect 3063 6452 3939 6472
rect 3063 6400 3467 6452
rect 3567 6400 3939 6452
rect 3063 6384 3939 6400
rect 3063 6343 3069 6384
rect 3023 6253 3069 6343
rect 3933 6343 3939 6384
rect 3973 6343 3979 6511
rect 3113 6325 3313 6335
rect 3101 6275 3113 6321
rect 3313 6315 3901 6321
rect 3889 6281 3901 6315
rect 3313 6275 3901 6281
rect 3113 6263 3313 6273
rect 3023 6085 3029 6253
rect 3063 6215 3069 6253
rect 3933 6253 3979 6343
rect 3933 6215 3939 6253
rect 3063 6200 3939 6215
rect 3063 6148 3464 6200
rect 3564 6185 3939 6200
rect 3973 6195 3979 6253
rect 3973 6185 3982 6195
rect 3564 6148 3930 6185
rect 3063 6127 3930 6148
rect 3063 6085 3069 6127
rect 3023 6073 3069 6085
rect 3465 6066 3565 6076
rect 3930 6075 3982 6085
rect 3933 6073 3979 6075
rect 3101 6057 3465 6063
rect 3565 6057 3901 6063
rect 3101 6023 3113 6057
rect 3889 6023 3901 6057
rect 3101 6017 3465 6023
rect 3565 6017 3901 6023
rect 3023 5995 3069 6007
rect 3465 6004 3565 6014
rect 3023 5827 3029 5995
rect 3063 5948 3069 5995
rect 3933 5995 3979 6007
rect 3933 5948 3939 5995
rect 3063 5860 3939 5948
rect 3063 5827 3069 5860
rect 3023 5737 3069 5827
rect 3933 5827 3939 5860
rect 3973 5827 3979 5995
rect 3689 5810 3889 5820
rect 3101 5799 3689 5805
rect 3101 5765 3113 5799
rect 3101 5759 3689 5765
rect 3889 5759 3901 5805
rect 3689 5744 3889 5754
rect 3023 5569 3029 5737
rect 3063 5704 3069 5737
rect 3933 5737 3979 5827
rect 3933 5704 3939 5737
rect 3063 5616 3939 5704
rect 3063 5569 3069 5616
rect 3023 5479 3069 5569
rect 3933 5569 3939 5616
rect 3973 5569 3979 5737
rect 3113 5556 3313 5566
rect 3101 5501 3113 5547
rect 3313 5541 3901 5547
rect 3889 5507 3901 5541
rect 3313 5501 3901 5507
rect 3113 5482 3313 5492
rect 3023 5311 3029 5479
rect 3063 5439 3069 5479
rect 3933 5479 3979 5569
rect 3933 5439 3939 5479
rect 3063 5351 3939 5439
rect 3063 5311 3069 5351
rect 3023 5221 3069 5311
rect 3933 5311 3939 5351
rect 3973 5311 3979 5479
rect 3689 5294 3889 5304
rect 3101 5283 3689 5289
rect 3101 5249 3113 5283
rect 3101 5243 3689 5249
rect 3889 5243 3901 5289
rect 3689 5228 3889 5238
rect 3023 5053 3029 5221
rect 3063 5188 3069 5221
rect 3933 5221 3979 5311
rect 3933 5188 3939 5221
rect 3063 5178 3939 5188
rect 3973 5184 3979 5221
rect 4156 5879 4208 6553
rect 3973 5178 3982 5184
rect 3063 5100 3930 5178
rect 3063 5053 3069 5100
rect 3023 5041 3069 5053
rect 3465 5034 3565 5044
rect 3930 5043 3982 5053
rect 4156 5105 4208 5779
rect 3933 5041 3979 5043
rect 3101 5025 3465 5031
rect 3565 5025 3901 5031
rect 3101 4991 3113 5025
rect 3889 4991 3901 5025
rect 3101 4985 3465 4991
rect 3565 4985 3901 4991
rect 3023 4963 3069 4975
rect 3465 4972 3565 4982
rect 3023 4795 3029 4963
rect 3063 4922 3069 4963
rect 3933 4963 3979 4975
rect 3933 4922 3939 4963
rect 3063 4909 3939 4922
rect 3063 4857 3462 4909
rect 3562 4857 3939 4909
rect 3063 4834 3939 4857
rect 3063 4795 3069 4834
rect 3023 4705 3069 4795
rect 3933 4795 3939 4834
rect 3973 4795 3979 4963
rect 3113 4776 3313 4786
rect 3101 4727 3113 4773
rect 3313 4767 3901 4773
rect 3889 4733 3901 4767
rect 3313 4727 3901 4733
rect 3113 4714 3313 4724
rect 3023 4537 3029 4705
rect 3063 4665 3069 4705
rect 3933 4705 3979 4795
rect 3933 4665 3939 4705
rect 3063 4647 3939 4665
rect 3063 4595 3459 4647
rect 3564 4637 3939 4647
rect 3973 4647 3979 4705
rect 3973 4637 3982 4647
rect 3564 4595 3930 4637
rect 3063 4577 3930 4595
rect 3063 4537 3069 4577
rect 3023 4525 3069 4537
rect 3465 4518 3565 4528
rect 3930 4527 3982 4537
rect 3933 4525 3979 4527
rect 3101 4509 3465 4515
rect 3565 4509 3901 4515
rect 3101 4475 3113 4509
rect 3889 4475 3901 4509
rect 3101 4469 3465 4475
rect 3565 4469 3901 4475
rect 3023 4447 3069 4459
rect 3465 4456 3565 4466
rect 3023 4279 3029 4447
rect 3063 4391 3069 4447
rect 3933 4447 3979 4459
rect 3933 4391 3939 4447
rect 3063 4303 3939 4391
rect 3063 4279 3069 4303
rect 3023 4189 3069 4279
rect 3933 4279 3939 4303
rect 3973 4279 3979 4447
rect 3689 4262 3889 4272
rect 3101 4251 3689 4257
rect 3101 4217 3113 4251
rect 3101 4211 3689 4217
rect 3889 4211 3901 4257
rect 3689 4196 3889 4206
rect 3023 4021 3029 4189
rect 3063 4148 3069 4189
rect 3933 4189 3979 4279
rect 3933 4148 3939 4189
rect 3063 4121 3939 4148
rect 3973 4131 3979 4189
rect 4156 4331 4208 5005
rect 3973 4121 3982 4131
rect 3063 4060 3930 4121
rect 3063 4021 3069 4060
rect 3023 4009 3069 4021
rect 3113 4008 3313 4018
rect 3930 4011 3982 4021
rect 4156 4073 4208 4231
rect 3933 4009 3979 4011
rect 3101 3953 3113 3999
rect 3313 3993 3901 3999
rect 3889 3959 3901 3993
rect 4156 3963 4208 3973
rect 4301 10007 4353 10129
rect 4504 10123 4550 10135
rect 5170 10132 5370 10142
rect 4504 10065 4510 10123
rect 4501 10055 4510 10065
rect 4544 10078 4550 10123
rect 5414 10123 5460 10135
rect 5414 10078 5420 10123
rect 4544 10059 5420 10078
rect 4544 10055 4897 10059
rect 4553 10007 4897 10055
rect 4997 10007 5420 10059
rect 4553 9990 5420 10007
rect 4501 9945 4553 9955
rect 5414 9955 5420 9990
rect 5454 9955 5460 10123
rect 4504 9943 4550 9945
rect 4895 9936 4995 9946
rect 5414 9943 5460 9955
rect 4301 9233 4353 9907
rect 4582 9927 4895 9933
rect 4995 9927 5382 9933
rect 4582 9893 4594 9927
rect 5370 9893 5382 9927
rect 4582 9887 4895 9893
rect 4995 9887 5382 9893
rect 4504 9865 4550 9877
rect 4895 9874 4995 9884
rect 4504 9697 4510 9865
rect 4544 9826 4550 9865
rect 5414 9865 5460 9877
rect 5414 9826 5420 9865
rect 4544 9738 5420 9826
rect 4544 9697 4550 9738
rect 4504 9607 4550 9697
rect 5414 9697 5420 9738
rect 5454 9697 5460 9865
rect 5169 9680 5369 9690
rect 4582 9669 5169 9675
rect 5369 9669 5382 9675
rect 4582 9635 4594 9669
rect 5370 9635 5382 9669
rect 4582 9629 5169 9635
rect 5369 9629 5382 9635
rect 5169 9614 5369 9624
rect 4504 9439 4510 9607
rect 4544 9577 4550 9607
rect 5414 9607 5460 9697
rect 5414 9577 5420 9607
rect 4544 9489 5420 9577
rect 4544 9439 4550 9489
rect 4504 9349 4550 9439
rect 5414 9439 5420 9489
rect 5454 9439 5460 9607
rect 4594 9426 4794 9436
rect 4582 9371 4594 9417
rect 4794 9411 5382 9417
rect 5370 9377 5382 9411
rect 4794 9371 5382 9377
rect 4594 9352 4794 9362
rect 4504 9181 4510 9349
rect 4544 9307 4550 9349
rect 5414 9349 5460 9439
rect 5414 9307 5420 9349
rect 4544 9219 5420 9307
rect 4544 9181 4550 9219
rect 4504 9133 4550 9181
rect 5414 9181 5420 9219
rect 5454 9181 5460 9349
rect 5170 9164 5370 9174
rect 4582 9153 5170 9159
rect 4301 8459 4353 9133
rect 4501 9123 4553 9133
rect 4582 9119 4594 9153
rect 4582 9113 5170 9119
rect 5370 9113 5382 9159
rect 5170 9098 5370 9108
rect 5414 9091 5460 9181
rect 5414 9058 5420 9091
rect 4553 8970 5420 9058
rect 4501 8913 4553 8923
rect 5414 8923 5420 8970
rect 5454 8923 5460 9091
rect 4504 8911 4550 8913
rect 4895 8904 4995 8914
rect 5414 8911 5460 8923
rect 4582 8895 4895 8901
rect 4995 8895 5382 8901
rect 4582 8861 4594 8895
rect 5370 8861 5382 8895
rect 4582 8855 4895 8861
rect 4995 8855 5382 8861
rect 4504 8833 4550 8845
rect 4895 8842 4995 8852
rect 4504 8665 4510 8833
rect 4544 8795 4550 8833
rect 5414 8833 5460 8845
rect 5414 8795 5420 8833
rect 4544 8781 5420 8795
rect 4544 8729 4894 8781
rect 4994 8729 5420 8781
rect 4544 8707 5420 8729
rect 4544 8665 4550 8707
rect 4504 8575 4550 8665
rect 5414 8665 5420 8707
rect 5454 8665 5460 8833
rect 5170 8646 5370 8656
rect 4582 8637 5170 8643
rect 4582 8603 4594 8637
rect 4582 8597 5170 8603
rect 5370 8597 5382 8643
rect 5170 8584 5370 8594
rect 4504 8517 4510 8575
rect 4501 8507 4510 8517
rect 4544 8541 4550 8575
rect 5414 8575 5460 8665
rect 5414 8541 5420 8575
rect 4544 8525 5420 8541
rect 4544 8507 4893 8525
rect 4553 8473 4893 8507
rect 4993 8473 5420 8525
rect 4553 8453 5420 8473
rect 4501 8397 4553 8407
rect 5414 8407 5420 8453
rect 5454 8407 5460 8575
rect 4504 8395 4550 8397
rect 4895 8388 4995 8398
rect 5414 8395 5460 8407
rect 4301 7685 4353 8359
rect 4582 8379 4895 8385
rect 4995 8379 5382 8385
rect 4582 8345 4594 8379
rect 5370 8345 5382 8379
rect 4582 8339 4895 8345
rect 4995 8339 5382 8345
rect 4301 6911 4353 7585
rect 4504 8317 4550 8329
rect 4895 8326 4995 8336
rect 4504 8149 4510 8317
rect 4544 8274 4550 8317
rect 5414 8317 5460 8329
rect 5414 8274 5420 8317
rect 4544 8186 5420 8274
rect 4544 8149 4550 8186
rect 4504 8059 4550 8149
rect 5414 8149 5420 8186
rect 5454 8149 5460 8317
rect 5170 8132 5370 8142
rect 4582 8121 5170 8127
rect 4582 8087 4594 8121
rect 4582 8081 5170 8087
rect 5370 8081 5382 8127
rect 5170 8066 5370 8076
rect 4504 7891 4510 8059
rect 4544 8021 4550 8059
rect 5414 8059 5460 8149
rect 5414 8021 5420 8059
rect 4544 7933 5420 8021
rect 4544 7891 4550 7933
rect 4504 7801 4550 7891
rect 5414 7891 5420 7933
rect 5454 7891 5460 8059
rect 4594 7878 4794 7888
rect 4582 7823 4594 7869
rect 4794 7863 5382 7869
rect 5370 7829 5382 7863
rect 4794 7823 5382 7829
rect 4594 7804 4794 7814
rect 4504 7633 4510 7801
rect 4544 7769 4550 7801
rect 5414 7801 5460 7891
rect 5414 7769 5420 7801
rect 4544 7681 5420 7769
rect 4544 7633 4550 7681
rect 4504 7569 4550 7633
rect 5414 7633 5420 7681
rect 5454 7633 5460 7801
rect 5170 7616 5370 7626
rect 4582 7605 5170 7611
rect 4582 7571 4594 7605
rect 4501 7559 4553 7569
rect 4582 7565 5170 7571
rect 5370 7565 5382 7611
rect 5170 7550 5370 7560
rect 5414 7543 5460 7633
rect 5414 7498 5420 7543
rect 4553 7410 5420 7498
rect 4501 7365 4553 7375
rect 5414 7375 5420 7410
rect 5454 7375 5460 7543
rect 4504 7363 4550 7365
rect 4895 7356 4995 7366
rect 5414 7363 5460 7375
rect 4582 7347 4895 7353
rect 4995 7347 5382 7353
rect 4582 7313 4594 7347
rect 5370 7313 5382 7347
rect 4582 7307 4895 7313
rect 4995 7307 5382 7313
rect 4504 7285 4550 7297
rect 4895 7294 4995 7304
rect 4504 7117 4510 7285
rect 4544 7252 4550 7285
rect 5414 7285 5460 7297
rect 5414 7252 5420 7285
rect 4544 7239 5420 7252
rect 4544 7187 4895 7239
rect 4995 7187 5420 7239
rect 4544 7171 5420 7187
rect 4544 7117 4550 7171
rect 4504 7027 4550 7117
rect 5414 7117 5420 7171
rect 5454 7117 5460 7285
rect 5170 7098 5370 7108
rect 4582 7089 5170 7095
rect 4582 7055 4594 7089
rect 4582 7049 5170 7055
rect 5370 7049 5382 7095
rect 5170 7036 5370 7046
rect 4504 6969 4510 7027
rect 4501 6959 4510 6969
rect 4544 6992 4550 7027
rect 5414 7027 5460 7117
rect 5414 6992 5420 7027
rect 4544 6977 5420 6992
rect 4544 6959 4897 6977
rect 4553 6925 4897 6959
rect 4997 6925 5420 6977
rect 4553 6911 5420 6925
rect 4501 6849 4553 6859
rect 5414 6859 5420 6911
rect 5454 6859 5460 7027
rect 4504 6847 4550 6849
rect 4894 6840 4994 6850
rect 5414 6847 5460 6859
rect 4301 6137 4353 6811
rect 4582 6831 4894 6837
rect 4994 6831 5382 6837
rect 4582 6797 4594 6831
rect 5370 6797 5382 6831
rect 4582 6791 4894 6797
rect 4994 6791 5382 6797
rect 4301 5363 4353 6037
rect 4504 6769 4550 6781
rect 4894 6778 4994 6788
rect 4504 6601 4510 6769
rect 4544 6730 4550 6769
rect 5414 6769 5460 6781
rect 5414 6730 5420 6769
rect 4544 6642 5420 6730
rect 4544 6601 4550 6642
rect 4504 6511 4550 6601
rect 5414 6601 5420 6642
rect 5454 6601 5460 6769
rect 5170 6584 5370 6594
rect 4582 6573 5170 6579
rect 4582 6539 4594 6573
rect 4582 6533 5170 6539
rect 5370 6533 5382 6579
rect 5170 6518 5370 6528
rect 4504 6343 4510 6511
rect 4544 6474 4550 6511
rect 5414 6511 5460 6601
rect 5414 6474 5420 6511
rect 4544 6386 5420 6474
rect 4544 6343 4550 6386
rect 4504 6253 4550 6343
rect 5414 6343 5420 6386
rect 5454 6343 5460 6511
rect 4594 6330 4794 6340
rect 4582 6275 4594 6321
rect 4794 6315 5382 6321
rect 5370 6281 5382 6315
rect 4794 6275 5382 6281
rect 4594 6256 4794 6266
rect 4504 6085 4510 6253
rect 4544 6213 4550 6253
rect 5414 6253 5460 6343
rect 5414 6213 5420 6253
rect 4544 6125 5420 6213
rect 4544 6085 4550 6125
rect 4504 6021 4550 6085
rect 5414 6085 5420 6125
rect 5454 6085 5460 6253
rect 5170 6068 5370 6078
rect 4582 6057 5170 6063
rect 4582 6023 4594 6057
rect 4501 6011 4553 6021
rect 4582 6017 5170 6023
rect 5370 6017 5382 6063
rect 5170 6002 5370 6012
rect 5414 5995 5460 6085
rect 5414 5958 5420 5995
rect 4553 5870 5420 5958
rect 4501 5817 4553 5827
rect 5414 5827 5420 5870
rect 5454 5827 5460 5995
rect 4504 5815 4550 5817
rect 4895 5808 4995 5818
rect 5414 5815 5460 5827
rect 4582 5799 4895 5805
rect 4995 5799 5382 5805
rect 4582 5765 4594 5799
rect 5370 5765 5382 5799
rect 4582 5759 4895 5765
rect 4995 5759 5382 5765
rect 4504 5737 4550 5749
rect 4895 5746 4995 5756
rect 4504 5569 4510 5737
rect 4544 5703 4550 5737
rect 5414 5737 5460 5749
rect 5414 5703 5420 5737
rect 4544 5681 5420 5703
rect 4544 5629 4897 5681
rect 4997 5629 5420 5681
rect 4544 5597 5420 5629
rect 4544 5569 4550 5597
rect 4504 5479 4550 5569
rect 5414 5569 5420 5597
rect 5454 5569 5460 5737
rect 5170 5550 5370 5560
rect 4582 5541 5170 5547
rect 4582 5507 4594 5541
rect 4582 5501 5170 5507
rect 5370 5501 5382 5547
rect 5170 5488 5370 5498
rect 4504 5421 4510 5479
rect 4501 5411 4510 5421
rect 4544 5448 4550 5479
rect 5414 5479 5460 5569
rect 5414 5448 5420 5479
rect 4544 5426 5420 5448
rect 4544 5411 4895 5426
rect 4553 5374 4895 5411
rect 4995 5374 5420 5426
rect 4553 5342 5420 5374
rect 4501 5301 4553 5311
rect 5414 5311 5420 5342
rect 5454 5311 5460 5479
rect 4504 5299 4550 5301
rect 4895 5292 4995 5302
rect 5414 5299 5460 5311
rect 4301 4589 4353 5263
rect 4582 5283 4895 5289
rect 4995 5283 5382 5289
rect 4582 5249 4594 5283
rect 5370 5249 5382 5283
rect 4582 5243 4895 5249
rect 4995 5243 5382 5249
rect 4301 4073 4353 4489
rect 4504 5221 4550 5233
rect 4895 5230 4995 5240
rect 4504 5053 4510 5221
rect 4544 5178 4550 5221
rect 5414 5221 5460 5233
rect 5414 5178 5420 5221
rect 4544 5090 5420 5178
rect 4544 5053 4550 5090
rect 4504 4963 4550 5053
rect 5414 5053 5420 5090
rect 5454 5053 5460 5221
rect 5170 5036 5370 5046
rect 4582 5025 5170 5031
rect 4582 4991 4594 5025
rect 4582 4985 5170 4991
rect 5370 4985 5382 5031
rect 5170 4970 5370 4980
rect 4504 4795 4510 4963
rect 4544 4922 4550 4963
rect 5414 4963 5460 5053
rect 5414 4922 5420 4963
rect 4544 4834 5420 4922
rect 4544 4795 4550 4834
rect 4504 4705 4550 4795
rect 5414 4795 5420 4834
rect 5454 4795 5460 4963
rect 4594 4782 4794 4792
rect 4582 4727 4594 4773
rect 4794 4767 5382 4773
rect 5370 4733 5382 4767
rect 4794 4727 5382 4733
rect 4594 4708 4794 4718
rect 4504 4537 4510 4705
rect 4544 4663 4550 4705
rect 5414 4705 5460 4795
rect 5414 4663 5420 4705
rect 4544 4575 5420 4663
rect 4544 4537 4550 4575
rect 4504 4473 4550 4537
rect 5414 4537 5420 4575
rect 5454 4537 5460 4705
rect 5170 4520 5370 4530
rect 4582 4509 5170 4515
rect 4582 4475 4594 4509
rect 4501 4463 4553 4473
rect 4582 4469 5170 4475
rect 5370 4469 5382 4515
rect 5170 4454 5370 4464
rect 5414 4447 5460 4537
rect 5414 4403 5420 4447
rect 4553 4315 5420 4403
rect 4501 4269 4553 4279
rect 5414 4279 5420 4315
rect 5454 4279 5460 4447
rect 4504 4267 4550 4269
rect 4895 4260 4995 4270
rect 5414 4267 5460 4279
rect 4582 4251 4895 4257
rect 4995 4251 5382 4257
rect 4582 4217 4594 4251
rect 5370 4217 5382 4251
rect 4582 4211 4895 4217
rect 4995 4211 5382 4217
rect 4504 4189 4550 4201
rect 4895 4198 4995 4208
rect 4504 4131 4510 4189
rect 4501 4121 4510 4131
rect 4544 4150 4550 4189
rect 5414 4189 5460 4201
rect 5414 4150 5420 4189
rect 4544 4134 5420 4150
rect 4544 4121 4893 4134
rect 4553 4082 4893 4121
rect 4993 4082 5420 4134
rect 4553 4062 5420 4082
rect 4501 4011 4553 4021
rect 5414 4021 5420 4062
rect 5454 4021 5460 4189
rect 4504 4009 4550 4011
rect 5170 4002 5370 4012
rect 5414 4009 5460 4021
rect 4301 3963 4353 3973
rect 4582 3993 5170 3999
rect 3313 3953 3901 3959
rect 4582 3959 4594 3993
rect 4582 3953 5170 3959
rect 3113 3934 3313 3944
rect 5370 3953 5382 3999
rect 5170 3940 5370 3950
rect 5623 3873 5629 10214
rect 5741 3873 5747 10214
rect 5784 10222 5892 10234
rect 5784 9695 5790 10222
rect 5886 9695 5892 10222
rect 5784 9683 5892 9695
rect 6210 10086 6262 10268
rect 6390 10248 6402 10368
rect 6881 10248 6893 10368
rect 7419 10303 7606 10309
rect 6390 10242 6893 10248
rect 6973 10271 7133 10283
rect 6402 10238 6881 10242
rect 6210 10055 6820 10086
rect 6210 10021 6255 10055
rect 6289 10021 6355 10055
rect 6389 10021 6455 10055
rect 6489 10021 6555 10055
rect 6589 10021 6655 10055
rect 6689 10021 6755 10055
rect 6789 10021 6820 10055
rect 6210 9955 6820 10021
rect 6210 9921 6255 9955
rect 6289 9921 6355 9955
rect 6389 9921 6455 9955
rect 6489 9921 6555 9955
rect 6589 9921 6655 9955
rect 6689 9921 6755 9955
rect 6789 9921 6820 9955
rect 6210 9855 6820 9921
rect 6210 9821 6255 9855
rect 6289 9821 6355 9855
rect 6389 9821 6455 9855
rect 6489 9821 6555 9855
rect 6589 9821 6655 9855
rect 6689 9821 6755 9855
rect 6789 9821 6820 9855
rect 6210 9755 6820 9821
rect 6210 9721 6255 9755
rect 6289 9721 6355 9755
rect 6389 9721 6455 9755
rect 6489 9721 6555 9755
rect 6589 9721 6655 9755
rect 6689 9721 6755 9755
rect 6789 9721 6820 9755
rect 6210 9655 6820 9721
rect 6210 9621 6255 9655
rect 6289 9621 6355 9655
rect 6389 9621 6455 9655
rect 6489 9621 6555 9655
rect 6589 9621 6655 9655
rect 6689 9621 6755 9655
rect 6789 9621 6820 9655
rect 6210 9588 6820 9621
rect 6210 9514 6215 9588
rect 6815 9514 6820 9588
rect 6210 9476 6820 9514
rect 6973 9446 6979 10271
rect 7127 9446 7133 10271
rect 7419 10269 7518 10303
rect 7594 10269 7606 10303
rect 7419 10263 7606 10269
rect 7419 10244 7465 10263
rect 7398 10241 7465 10244
rect 7398 10234 7425 10241
rect 7459 10234 7465 10241
rect 7463 10194 7465 10234
rect 7647 10241 7693 10253
rect 7647 10194 7653 10241
rect 7463 9912 7653 10194
rect 7463 9875 7465 9912
rect 7398 9873 7425 9875
rect 7459 9873 7465 9875
rect 7398 9865 7465 9873
rect 7419 9790 7465 9865
rect 7647 9873 7653 9912
rect 7687 9873 7693 10241
rect 7518 9854 7594 9864
rect 7647 9861 7693 9873
rect 7506 9805 7518 9851
rect 7594 9805 7606 9851
rect 7518 9792 7594 9802
rect 6973 9434 7133 9446
rect 7398 9783 7465 9790
rect 7398 9780 7425 9783
rect 7459 9780 7465 9783
rect 7463 9747 7465 9780
rect 7647 9783 7693 9795
rect 7647 9747 7653 9783
rect 7463 9465 7653 9747
rect 7463 9421 7465 9465
rect 7398 9415 7425 9421
rect 7459 9415 7465 9421
rect 7398 9411 7465 9415
rect 7419 9393 7465 9411
rect 7647 9415 7653 9465
rect 7687 9415 7693 9783
rect 7847 9499 7853 10480
rect 7647 9403 7693 9415
rect 7845 9487 7853 9499
rect 7985 9499 7991 10480
rect 8058 10479 8218 10491
rect 7985 9487 7992 9499
rect 7419 9387 7606 9393
rect 7419 9353 7518 9387
rect 7594 9353 7606 9387
rect 7419 9347 7606 9353
rect 5969 9327 7012 9331
rect 5957 9321 7024 9327
rect 5957 9213 5969 9321
rect 7012 9213 7024 9321
rect 5957 9207 7024 9213
rect 5969 9203 7012 9207
rect 7419 9116 7465 9347
rect 7518 9193 7658 9203
rect 7506 9138 7518 9184
rect 7658 9178 7706 9184
rect 7694 9144 7706 9178
rect 7658 9138 7706 9144
rect 7518 9119 7658 9129
rect 7419 8948 7425 9116
rect 7459 9085 7465 9116
rect 7747 9116 7793 9128
rect 7747 9085 7753 9116
rect 7459 8967 7753 9085
rect 7459 8948 7465 8967
rect 7419 8858 7465 8948
rect 7747 8948 7753 8967
rect 7787 8948 7793 9116
rect 7554 8929 7694 8939
rect 7747 8936 7793 8948
rect 7506 8920 7554 8926
rect 7506 8886 7518 8920
rect 7506 8880 7554 8886
rect 7694 8880 7706 8926
rect 7554 8867 7694 8877
rect 7419 8690 7425 8858
rect 7459 8833 7465 8858
rect 7747 8858 7793 8870
rect 7747 8833 7753 8858
rect 7459 8715 7753 8833
rect 7459 8690 7465 8715
rect 5623 3861 5747 3873
rect 6365 8370 6568 8382
rect 2682 3817 2868 3829
rect 6365 2963 6371 8370
rect 6562 2963 6568 8370
rect 6731 8258 6791 8268
rect 6719 8209 6731 8255
rect 6791 8249 6919 8255
rect 6907 8215 6919 8249
rect 6791 8209 6919 8215
rect 6641 8187 6687 8199
rect 6731 8196 6791 8206
rect 6641 8019 6647 8187
rect 6681 8138 6687 8187
rect 6951 8187 6997 8199
rect 6951 8138 6957 8187
rect 6681 8071 6957 8138
rect 6681 8019 6687 8071
rect 6641 7929 6687 8019
rect 6951 8019 6957 8071
rect 6991 8019 6997 8187
rect 6731 8000 6791 8010
rect 6719 7951 6731 7997
rect 6791 7991 6919 7997
rect 6907 7957 6919 7991
rect 6791 7951 6919 7957
rect 6731 7938 6791 7948
rect 6641 7761 6647 7929
rect 6681 7880 6687 7929
rect 6951 7929 6997 8019
rect 6951 7880 6957 7929
rect 6681 7813 6957 7880
rect 6681 7761 6687 7813
rect 6641 7739 6687 7761
rect 6951 7761 6957 7813
rect 6991 7761 6997 7929
rect 6951 7752 6997 7761
rect 6847 7742 6997 7752
rect 6641 7733 6847 7739
rect 6641 7699 6731 7733
rect 6641 7693 6847 7699
rect 6641 7671 6687 7693
rect 6907 7690 6997 7742
rect 6847 7680 6997 7690
rect 6641 7503 6647 7671
rect 6681 7618 6687 7671
rect 6951 7671 6997 7680
rect 6951 7618 6957 7671
rect 6681 7551 6957 7618
rect 6681 7503 6687 7551
rect 6641 7413 6687 7503
rect 6951 7503 6957 7551
rect 6991 7503 6997 7671
rect 6731 7484 6791 7494
rect 6719 7435 6731 7481
rect 6791 7475 6919 7481
rect 6907 7441 6919 7475
rect 6791 7435 6919 7441
rect 6731 7422 6791 7432
rect 6641 7245 6647 7413
rect 6681 7361 6687 7413
rect 6951 7413 6997 7503
rect 6951 7361 6957 7413
rect 6681 7294 6957 7361
rect 6681 7245 6687 7294
rect 6641 7223 6687 7245
rect 6951 7245 6957 7294
rect 6991 7245 6997 7413
rect 6951 7236 6997 7245
rect 6847 7226 6997 7236
rect 6641 7217 6847 7223
rect 6641 7183 6731 7217
rect 6641 7177 6847 7183
rect 6641 7155 6687 7177
rect 6907 7174 6997 7226
rect 6847 7164 6997 7174
rect 6641 6987 6647 7155
rect 6681 7101 6687 7155
rect 6951 7155 6997 7164
rect 6951 7101 6957 7155
rect 6681 7034 6957 7101
rect 6681 6987 6687 7034
rect 6641 6975 6687 6987
rect 6951 6987 6957 7034
rect 6991 6987 6997 7155
rect 6731 6968 6791 6978
rect 6951 6975 6997 6987
rect 7419 7871 7465 8690
rect 7747 8690 7753 8715
rect 7787 8690 7793 8858
rect 7518 8677 7658 8687
rect 7747 8678 7793 8690
rect 7506 8622 7518 8668
rect 7658 8662 7706 8668
rect 7694 8628 7706 8662
rect 7658 8622 7706 8628
rect 7518 8603 7658 8613
rect 7845 8501 7851 9487
rect 7986 8501 7992 9487
rect 7845 8489 7992 8501
rect 8058 8500 8064 10479
rect 8212 8500 8218 10479
rect 18028 10318 18175 10654
rect 18209 10318 18228 10654
rect 18028 10305 18228 10318
rect 18028 9274 18114 10305
rect 18405 10265 21644 10707
rect 21827 10654 21873 10666
rect 21813 10318 21823 10654
rect 21877 10318 21887 10654
rect 21827 10306 21873 10318
rect 22067 10265 25306 10707
rect 25471 10654 25673 10667
rect 25471 10318 25491 10654
rect 25525 10318 25673 10654
rect 25471 10307 25673 10318
rect 25485 10306 25531 10307
rect 18225 10259 21817 10265
rect 18225 10225 18237 10259
rect 21805 10225 21817 10259
rect 18225 10219 21817 10225
rect 21883 10259 25475 10265
rect 21883 10225 21895 10259
rect 25463 10225 25475 10259
rect 21883 10219 25475 10225
rect 18142 10166 18228 10178
rect 18142 10135 18175 10166
rect 18209 10135 18228 10166
rect 18218 9830 18228 10135
rect 18142 9817 18228 9830
rect 18405 9777 21644 10219
rect 21827 10166 21873 10178
rect 21813 9830 21823 10166
rect 21877 9830 21887 10166
rect 21827 9818 21873 9830
rect 22067 9777 25306 10219
rect 25473 10166 25559 10178
rect 25473 10125 25491 10166
rect 25525 10125 25559 10166
rect 25473 9830 25483 10125
rect 25473 9777 25559 9830
rect 18225 9771 25559 9777
rect 18225 9737 18237 9771
rect 21805 9737 21895 9771
rect 25463 9737 25559 9771
rect 18225 9731 25559 9737
rect 25587 9459 25673 10307
rect 18142 9458 25901 9459
rect 26488 9458 26498 9459
rect 18142 9452 26498 9458
rect 18451 9444 26498 9452
rect 18451 9377 18950 9444
rect 19299 9441 26498 9444
rect 19299 9377 24014 9441
rect 18451 9374 24014 9377
rect 24363 9374 26498 9441
rect 18451 9368 26498 9374
rect 18142 9359 26498 9368
rect 25886 9358 26498 9359
rect 26488 9298 26498 9358
rect 26678 9298 26688 9459
rect 18028 9258 25569 9274
rect 18028 9254 24434 9258
rect 18028 9187 19377 9254
rect 19726 9191 24434 9254
rect 24783 9191 25148 9258
rect 19726 9188 25148 9191
rect 25538 9188 25569 9258
rect 19726 9187 25569 9188
rect 18028 9174 25569 9187
rect 19435 8866 21827 8872
rect 19435 8832 19447 8866
rect 21815 8832 21827 8866
rect 19435 8826 21827 8832
rect 21893 8866 24285 8872
rect 21893 8832 21905 8866
rect 24273 8832 24285 8866
rect 21893 8826 24285 8832
rect 19379 8782 19425 8794
rect 8058 8488 8218 8500
rect 19331 8214 19341 8782
rect 19427 8214 19437 8782
rect 7571 7942 7694 7952
rect 7506 7933 7571 7939
rect 7959 7940 8110 7952
rect 7506 7899 7518 7933
rect 7506 7893 7571 7899
rect 7694 7893 7706 7939
rect 7571 7880 7694 7890
rect 7419 7503 7425 7871
rect 7459 7833 7465 7871
rect 7747 7871 7793 7883
rect 7747 7833 7753 7871
rect 7459 7554 7753 7833
rect 7459 7503 7465 7554
rect 6719 6919 6731 6965
rect 6791 6959 6919 6965
rect 6907 6925 6919 6959
rect 6791 6919 6919 6925
rect 6641 6897 6687 6909
rect 6731 6906 6791 6916
rect 6641 6729 6647 6897
rect 6681 6849 6687 6897
rect 6951 6897 6997 6909
rect 6951 6849 6957 6897
rect 6681 6782 6957 6849
rect 6681 6729 6687 6782
rect 6641 6639 6687 6729
rect 6951 6729 6957 6782
rect 6991 6729 6997 6897
rect 6731 6710 6791 6720
rect 6719 6661 6731 6707
rect 6791 6701 6919 6707
rect 6907 6667 6919 6701
rect 6791 6661 6919 6667
rect 6731 6648 6791 6658
rect 6641 6471 6647 6639
rect 6681 6595 6687 6639
rect 6951 6639 6997 6729
rect 6951 6595 6957 6639
rect 6681 6528 6957 6595
rect 6681 6471 6687 6528
rect 6641 6449 6687 6471
rect 6951 6471 6957 6528
rect 6991 6471 6997 6639
rect 6951 6462 6997 6471
rect 6847 6452 6997 6462
rect 6641 6443 6847 6449
rect 6641 6409 6731 6443
rect 6641 6403 6847 6409
rect 6641 6381 6687 6403
rect 6907 6400 6997 6452
rect 6847 6390 6997 6400
rect 6641 6213 6647 6381
rect 6681 6334 6687 6381
rect 6951 6381 6997 6390
rect 6951 6334 6957 6381
rect 6681 6267 6957 6334
rect 6681 6213 6687 6267
rect 6641 6123 6687 6213
rect 6951 6213 6957 6267
rect 6991 6213 6997 6381
rect 6731 6194 6791 6204
rect 6719 6145 6731 6191
rect 6791 6185 6919 6191
rect 6907 6151 6919 6185
rect 6791 6145 6919 6151
rect 6731 6132 6791 6142
rect 6641 5955 6647 6123
rect 6681 6081 6687 6123
rect 6951 6123 6997 6213
rect 6951 6081 6957 6123
rect 6681 6014 6957 6081
rect 6681 5955 6687 6014
rect 6641 5933 6687 5955
rect 6951 5955 6957 6014
rect 6991 5955 6997 6123
rect 6951 5946 6997 5955
rect 6847 5936 6997 5946
rect 6641 5927 6847 5933
rect 6641 5893 6731 5927
rect 6641 5887 6847 5893
rect 6641 5865 6687 5887
rect 6907 5884 6997 5936
rect 6847 5874 6997 5884
rect 6641 5697 6647 5865
rect 6681 5819 6687 5865
rect 6951 5865 6997 5874
rect 6951 5819 6957 5865
rect 6681 5752 6957 5819
rect 6681 5697 6687 5752
rect 6641 5685 6687 5697
rect 6951 5697 6957 5752
rect 6991 5697 6997 5865
rect 6731 5678 6791 5688
rect 6951 5685 6997 5697
rect 7419 6581 7465 7503
rect 7747 7503 7753 7554
rect 7787 7503 7793 7871
rect 7518 7484 7631 7494
rect 7747 7491 7793 7503
rect 7506 7435 7518 7481
rect 7631 7475 7706 7481
rect 7694 7441 7706 7475
rect 7631 7435 7706 7441
rect 7518 7422 7631 7432
rect 7571 6652 7694 6662
rect 7506 6643 7571 6649
rect 7506 6609 7518 6643
rect 7506 6603 7571 6609
rect 7694 6603 7706 6649
rect 7571 6590 7694 6600
rect 7419 6213 7425 6581
rect 7459 6535 7465 6581
rect 7747 6581 7793 6593
rect 7747 6535 7753 6581
rect 7459 6256 7753 6535
rect 7459 6213 7465 6256
rect 6719 5629 6731 5675
rect 6791 5669 6919 5675
rect 6907 5635 6919 5669
rect 6791 5629 6919 5635
rect 6641 5607 6687 5619
rect 6731 5616 6791 5626
rect 6641 5439 6647 5607
rect 6681 5561 6687 5607
rect 6951 5607 6997 5619
rect 6951 5561 6957 5607
rect 6681 5494 6957 5561
rect 6681 5439 6687 5494
rect 6641 5349 6687 5439
rect 6951 5439 6957 5494
rect 6991 5439 6997 5607
rect 6731 5420 6791 5430
rect 6719 5371 6731 5417
rect 6791 5411 6919 5417
rect 6907 5377 6919 5411
rect 6791 5371 6919 5377
rect 6731 5358 6791 5368
rect 6641 5181 6647 5349
rect 6681 5304 6687 5349
rect 6951 5349 6997 5439
rect 6951 5304 6957 5349
rect 6681 5237 6957 5304
rect 6681 5181 6687 5237
rect 6641 5159 6687 5181
rect 6951 5181 6957 5237
rect 6991 5181 6997 5349
rect 6951 5172 6997 5181
rect 6847 5162 6997 5172
rect 6641 5153 6847 5159
rect 6641 5119 6731 5153
rect 6641 5113 6847 5119
rect 6641 5091 6687 5113
rect 6907 5110 6997 5162
rect 6847 5100 6997 5110
rect 6641 4923 6647 5091
rect 6681 5043 6687 5091
rect 6951 5091 6997 5100
rect 6951 5043 6957 5091
rect 6681 4976 6957 5043
rect 6681 4923 6687 4976
rect 6641 4833 6687 4923
rect 6951 4923 6957 4976
rect 6991 4923 6997 5091
rect 6731 4904 6791 4914
rect 6719 4855 6731 4901
rect 6791 4895 6919 4901
rect 6907 4861 6919 4895
rect 6791 4855 6919 4861
rect 6731 4842 6791 4852
rect 6641 4665 6647 4833
rect 6681 4784 6687 4833
rect 6951 4833 6997 4923
rect 6951 4784 6957 4833
rect 6681 4717 6957 4784
rect 6681 4665 6687 4717
rect 6641 4643 6687 4665
rect 6951 4665 6957 4717
rect 6991 4665 6997 4833
rect 6951 4656 6997 4665
rect 6847 4646 6997 4656
rect 6641 4637 6847 4643
rect 6641 4603 6731 4637
rect 6641 4597 6847 4603
rect 6641 4575 6687 4597
rect 6907 4594 6997 4646
rect 6847 4584 6997 4594
rect 6641 4407 6647 4575
rect 6681 4534 6687 4575
rect 6951 4575 6997 4584
rect 6951 4534 6957 4575
rect 6681 4467 6957 4534
rect 6681 4407 6687 4467
rect 6641 4395 6687 4407
rect 6951 4407 6957 4467
rect 6991 4407 6997 4575
rect 6731 4388 6791 4398
rect 6951 4395 6997 4407
rect 7419 5291 7465 6213
rect 7747 6213 7753 6256
rect 7787 6213 7793 6581
rect 7518 6194 7631 6204
rect 7747 6201 7793 6213
rect 7506 6145 7518 6191
rect 7631 6185 7706 6191
rect 7694 6151 7706 6185
rect 7631 6145 7706 6151
rect 7518 6132 7631 6142
rect 7571 5362 7694 5372
rect 7506 5353 7571 5359
rect 7506 5319 7518 5353
rect 7506 5313 7571 5319
rect 7694 5313 7706 5359
rect 7571 5300 7694 5310
rect 7419 4923 7425 5291
rect 7459 5254 7465 5291
rect 7747 5291 7793 5303
rect 7747 5254 7753 5291
rect 7459 4975 7753 5254
rect 7459 4923 7465 4975
rect 6719 4339 6731 4385
rect 6791 4379 6919 4385
rect 6907 4345 6919 4379
rect 6791 4339 6919 4345
rect 6641 4317 6687 4329
rect 6731 4326 6791 4336
rect 6641 4149 6647 4317
rect 6681 4274 6687 4317
rect 6951 4317 6997 4329
rect 6951 4274 6957 4317
rect 6681 4207 6957 4274
rect 6681 4149 6687 4207
rect 6641 4059 6687 4149
rect 6951 4149 6957 4207
rect 6991 4149 6997 4317
rect 6731 4130 6791 4140
rect 6719 4081 6731 4127
rect 6791 4121 6919 4127
rect 6907 4087 6919 4121
rect 6791 4081 6919 4087
rect 6731 4068 6791 4078
rect 6641 3891 6647 4059
rect 6681 4012 6687 4059
rect 6951 4059 6997 4149
rect 6951 4012 6957 4059
rect 6681 3945 6957 4012
rect 6681 3891 6687 3945
rect 6641 3869 6687 3891
rect 6951 3891 6957 3945
rect 6991 3891 6997 4059
rect 6951 3882 6997 3891
rect 6847 3872 6997 3882
rect 6641 3863 6847 3869
rect 6641 3829 6731 3863
rect 6641 3823 6847 3829
rect 6641 3801 6687 3823
rect 6907 3820 6997 3872
rect 6847 3810 6997 3820
rect 6641 3633 6647 3801
rect 6681 3752 6687 3801
rect 6951 3801 6997 3810
rect 6951 3752 6957 3801
rect 6681 3685 6957 3752
rect 6681 3633 6687 3685
rect 6641 3543 6687 3633
rect 6951 3633 6957 3685
rect 6991 3633 6997 3801
rect 6731 3614 6791 3624
rect 6719 3565 6731 3611
rect 6791 3605 6919 3611
rect 6907 3571 6919 3605
rect 6791 3565 6919 3571
rect 6731 3552 6791 3562
rect 6641 3375 6647 3543
rect 6681 3493 6687 3543
rect 6951 3543 6997 3633
rect 6951 3493 6957 3543
rect 6681 3426 6957 3493
rect 6681 3375 6687 3426
rect 6641 3353 6687 3375
rect 6951 3375 6957 3426
rect 6991 3375 6997 3543
rect 6951 3366 6997 3375
rect 6847 3356 6997 3366
rect 6641 3347 6847 3353
rect 6641 3313 6731 3347
rect 6641 3307 6847 3313
rect 6641 3285 6687 3307
rect 6907 3304 6997 3356
rect 6847 3294 6997 3304
rect 6641 3117 6647 3285
rect 6681 3226 6687 3285
rect 6951 3285 6997 3294
rect 6951 3226 6957 3285
rect 6681 3159 6957 3226
rect 6681 3117 6687 3159
rect 6641 3105 6687 3117
rect 6951 3117 6957 3159
rect 6991 3117 6997 3285
rect 6731 3098 6791 3108
rect 6719 3049 6731 3095
rect 6847 3098 6907 3108
rect 6951 3105 6997 3117
rect 7419 4001 7465 4923
rect 7747 4923 7753 4975
rect 7787 4923 7793 5291
rect 7518 4904 7631 4914
rect 7747 4911 7793 4923
rect 7506 4855 7518 4901
rect 7631 4895 7706 4901
rect 7694 4861 7706 4895
rect 7631 4855 7706 4861
rect 7518 4842 7631 4852
rect 7959 4287 7965 7940
rect 7955 4202 7959 4260
rect 7570 4072 7694 4082
rect 7506 4063 7570 4069
rect 7506 4029 7518 4063
rect 7506 4023 7570 4029
rect 7694 4023 7706 4069
rect 7570 4010 7694 4020
rect 7419 3633 7425 4001
rect 7459 3944 7465 4001
rect 7747 4001 7793 4013
rect 7747 3944 7753 4001
rect 7459 3665 7753 3944
rect 7459 3633 7465 3665
rect 7419 3420 7465 3633
rect 7747 3633 7753 3665
rect 7787 3633 7793 4001
rect 7518 3614 7641 3624
rect 7747 3621 7793 3633
rect 7506 3565 7518 3611
rect 7641 3605 7706 3611
rect 7694 3571 7706 3605
rect 7641 3565 7706 3571
rect 7518 3552 7641 3562
rect 7571 3491 7694 3501
rect 7506 3482 7571 3488
rect 7506 3448 7518 3482
rect 7506 3442 7571 3448
rect 7694 3442 7706 3488
rect 7571 3429 7694 3439
rect 6791 3089 6847 3095
rect 6791 3049 6847 3055
rect 6731 3036 6791 3046
rect 6907 3049 6919 3095
rect 7419 3052 7425 3420
rect 7459 3368 7465 3420
rect 7747 3420 7793 3432
rect 7747 3368 7753 3420
rect 7459 3089 7753 3368
rect 7459 3052 7465 3089
rect 6847 3036 6907 3046
rect 7419 3035 7465 3052
rect 7747 3052 7753 3089
rect 7787 3052 7793 3420
rect 7518 3033 7641 3043
rect 7747 3040 7793 3052
rect 7506 2984 7518 3030
rect 7641 3024 7706 3030
rect 7694 2990 7706 3024
rect 7641 2984 7706 2990
rect 7518 2971 7641 2981
rect 6365 2951 6568 2963
rect 8104 4287 8110 7940
rect 19331 7648 19385 8214
rect 19379 7606 19385 7648
rect 19419 7648 19437 8214
rect 19419 7606 19425 7648
rect 19379 7594 19425 7606
rect 20083 7568 21168 8826
rect 21837 8782 21883 8794
rect 21837 7957 21843 8782
rect 21877 7957 21883 8782
rect 21825 7638 21835 7957
rect 21887 7638 21897 7957
rect 21837 7606 21843 7638
rect 21877 7606 21883 7638
rect 21837 7594 21883 7606
rect 22587 7568 23674 8826
rect 24295 8782 24341 8794
rect 24283 8214 24293 8782
rect 24379 8214 24389 8782
rect 24283 7661 24301 8214
rect 24295 7606 24301 7661
rect 24335 7661 24389 8214
rect 24335 7606 24341 7661
rect 24295 7594 24341 7606
rect 19441 7562 19451 7568
rect 19435 7556 19451 7562
rect 19661 7562 21825 7568
rect 21895 7562 24063 7568
rect 19661 7556 21827 7562
rect 19435 7522 19447 7556
rect 21815 7522 21827 7556
rect 19435 7516 19451 7522
rect 19441 7511 19451 7516
rect 19661 7516 21827 7522
rect 21893 7556 24063 7562
rect 24273 7562 24283 7568
rect 21893 7522 21905 7556
rect 21893 7516 24063 7522
rect 19661 7511 21825 7516
rect 21895 7511 24063 7516
rect 24273 7516 24285 7562
rect 24273 7511 24283 7516
rect 19451 7450 21904 7454
rect 19451 7393 19474 7450
rect 19661 7393 21904 7450
rect 19451 7390 21904 7393
rect 22105 7390 22114 7454
rect 19451 7375 22114 7390
rect 18048 7275 18058 7286
rect 18046 7231 18058 7275
rect 18634 7275 18644 7286
rect 18634 7231 18646 7275
rect 18046 7229 18646 7231
rect 17968 7207 18014 7219
rect 17968 6239 17974 7207
rect 18008 7020 18014 7207
rect 18678 7207 18737 7219
rect 18678 7038 18684 7207
rect 18718 7038 18737 7207
rect 21604 7137 24273 7157
rect 21604 7135 24063 7137
rect 21814 7080 24063 7135
rect 21814 7078 24273 7080
rect 21604 7068 24273 7078
rect 18666 7020 18676 7038
rect 18008 6423 18676 7020
rect 18008 6239 18014 6423
rect 18666 6239 18676 6423
rect 18728 6239 18738 7038
rect 19436 6997 21604 7003
rect 19434 6991 21604 6997
rect 21814 6997 21824 7003
rect 21894 6997 21904 7002
rect 19434 6957 19446 6991
rect 19434 6951 21604 6957
rect 19436 6946 21604 6951
rect 21814 6951 21826 6997
rect 21892 6951 21904 6997
rect 22114 6997 24282 7002
rect 22114 6991 24284 6997
rect 24272 6957 24284 6991
rect 21814 6946 21824 6951
rect 19378 6907 19424 6919
rect 17968 6227 18014 6239
rect 18678 6227 18737 6239
rect 18046 6211 18646 6217
rect 18046 6177 18058 6211
rect 18634 6177 18646 6211
rect 18046 6171 18646 6177
rect 19225 5835 19274 6907
rect 19426 5835 19436 6907
rect 19225 5766 19384 5835
rect 19378 5731 19384 5766
rect 19418 5766 19436 5835
rect 19418 5731 19424 5766
rect 19378 5719 19424 5731
rect 20078 5688 21165 6946
rect 21894 6945 21904 6951
rect 22114 6951 24284 6957
rect 22114 6945 24282 6951
rect 21836 6907 21882 6919
rect 21836 6876 21842 6907
rect 21876 6876 21882 6907
rect 21824 6557 21834 6876
rect 21886 6557 21896 6876
rect 21836 5731 21842 6557
rect 21876 5731 21882 6557
rect 21836 5719 21882 5731
rect 17820 5667 18397 5673
rect 17820 5573 17832 5667
rect 18385 5573 18397 5667
rect 19434 5636 19446 5688
rect 19926 5681 21826 5688
rect 21894 5687 21904 5689
rect 21814 5647 21826 5681
rect 19926 5636 21826 5647
rect 21892 5641 21904 5687
rect 22384 5687 22394 5689
rect 22578 5687 23665 6945
rect 24294 6907 24340 6919
rect 24281 5835 24291 6907
rect 24443 5835 24453 6907
rect 24294 5731 24300 5835
rect 24334 5731 24340 5835
rect 24294 5719 24340 5731
rect 22384 5681 24284 5687
rect 24272 5647 24284 5681
rect 21894 5637 21904 5641
rect 22384 5641 24284 5647
rect 22384 5637 22394 5641
rect 17820 5567 18397 5573
rect 17822 5432 24780 5438
rect 17822 5343 17834 5432
rect 24768 5343 24780 5432
rect 17822 5337 24780 5343
rect 8110 4202 8114 4260
rect 7959 2923 8110 2933
<< via1 >>
rect 11800 32809 14392 33012
rect 3401 30801 11199 30890
rect 7314 30104 7324 30440
rect 7324 30104 7358 30440
rect 7358 30104 7368 30440
rect 3633 29616 3666 29921
rect 3666 29616 3700 29921
rect 3700 29616 3709 29921
rect 7314 29616 7324 29952
rect 7324 29616 7358 29952
rect 7358 29616 7368 29952
rect 10974 29616 10982 29911
rect 10982 29616 11016 29911
rect 11016 29616 11050 29911
rect 11800 29401 11965 32809
rect 12122 29540 12138 30540
rect 12138 29540 12172 30540
rect 12172 29540 12186 30540
rect 12557 31916 12576 32516
rect 12576 31916 12610 32516
rect 12610 31916 12629 32516
rect 12999 30777 13014 31777
rect 13014 30777 13048 31777
rect 13048 30777 13063 31777
rect 13433 31916 13452 32516
rect 13452 31916 13486 32516
rect 13486 31916 13505 32516
rect 13875 29540 13890 30540
rect 13890 29540 13924 30540
rect 13924 29540 13939 30540
rect 12200 29481 12480 29490
rect 12200 29447 12480 29481
rect 12200 29438 12480 29447
rect 12638 29481 12918 29490
rect 12638 29447 12918 29481
rect 12638 29438 12918 29447
rect 13076 29481 13356 29490
rect 13076 29447 13356 29481
rect 13076 29438 13356 29447
rect 13514 29481 13794 29490
rect 13514 29447 13794 29481
rect 13514 29438 13794 29447
rect 3633 29154 3942 29238
rect 4441 29163 4790 29230
rect 9505 29160 9854 29227
rect 12200 29145 12300 29245
rect 12886 29145 12986 29245
rect 13324 29145 13424 29245
rect 13514 29145 13614 29245
rect 15339 29145 15621 29245
rect 4868 28973 5217 29040
rect 9925 28977 10274 29044
rect 10639 28974 11029 29044
rect 12448 28836 12548 28936
rect 12638 28836 12738 28936
rect 13076 28836 13176 28936
rect 13762 28836 13862 28936
rect 12268 28632 12548 28641
rect 4832 28000 4876 28568
rect 4876 28000 4910 28568
rect 4910 28000 4918 28568
rect 7326 27424 7334 27743
rect 7334 27424 7368 27743
rect 7368 27424 7378 27743
rect 12268 28598 12548 28632
rect 12268 28589 12548 28598
rect 12706 28632 12986 28641
rect 12706 28598 12986 28632
rect 12706 28589 12986 28598
rect 13144 28632 13424 28641
rect 13144 28598 13424 28632
rect 13144 28589 13424 28598
rect 13582 28632 13862 28641
rect 13582 28598 13862 28632
rect 13582 28589 13862 28598
rect 9784 28000 9792 28568
rect 9792 28000 9826 28568
rect 9826 28000 9870 28568
rect 4942 27342 5152 27354
rect 4942 27308 5152 27342
rect 4942 27297 5152 27308
rect 9554 27342 9764 27354
rect 9554 27308 9764 27342
rect 9554 27297 9764 27308
rect 4965 27179 5152 27236
rect 7395 27176 7596 27240
rect 3549 27055 4125 27072
rect 3549 27021 4125 27055
rect 3549 27017 4125 27021
rect 7095 26864 7305 26921
rect 9554 26866 9764 26923
rect 4167 26025 4175 26824
rect 4175 26025 4209 26824
rect 4209 26025 4219 26824
rect 7095 26777 7305 26789
rect 7095 26743 7305 26777
rect 7095 26732 7305 26743
rect 7395 26777 7605 26788
rect 7395 26743 7605 26777
rect 4765 25621 4875 26693
rect 4875 25621 4909 26693
rect 4909 25621 4917 26693
rect 7395 26731 7605 26743
rect 7325 26343 7333 26662
rect 7333 26343 7367 26662
rect 7367 26343 7377 26662
rect 3323 25359 3876 25453
rect 4937 25467 5417 25474
rect 4937 25433 5417 25467
rect 4937 25422 5417 25433
rect 7395 25467 7875 25475
rect 9782 25621 9791 26693
rect 9791 25621 9825 26693
rect 9825 25621 9934 26693
rect 7395 25433 7875 25467
rect 7395 25423 7875 25433
rect 11817 25407 11965 28583
rect 11816 25374 11965 25407
rect 12123 27539 12138 28539
rect 12138 27539 12172 28539
rect 12172 27539 12187 28539
rect 12557 25563 12576 26163
rect 12576 25563 12610 26163
rect 12610 25563 12629 26163
rect 12999 26379 13014 27379
rect 13014 26379 13048 27379
rect 13048 26379 13063 27379
rect 13432 25563 13452 26163
rect 13452 25563 13486 26163
rect 13486 25563 13504 26163
rect 13875 27539 13890 28539
rect 13890 27539 13924 28539
rect 13924 27539 13939 28539
rect 25403 28157 25662 28158
rect 20700 27793 25662 28157
rect 20700 27792 25504 27793
rect 15475 27207 19138 27498
rect 11816 25231 14381 25374
rect 11929 25230 14381 25231
rect 3325 25129 10259 25218
rect 16958 25985 16967 26985
rect 16967 25985 17001 26985
rect 17001 25985 17010 26985
rect 17376 25609 17385 26609
rect 17385 25609 17419 26609
rect 17419 25609 17428 26609
rect 17794 25985 17803 26985
rect 17803 25985 17837 26985
rect 17837 25985 17846 26985
rect 18212 25609 18221 26609
rect 18221 25609 18255 26609
rect 18255 25609 18264 26609
rect 18630 25985 18639 26985
rect 18639 25985 18673 26985
rect 18673 25985 18682 26985
rect 18851 25691 19138 27207
rect 18838 25506 18962 25565
rect 20762 25590 20879 27792
rect 21045 27054 21060 27254
rect 21060 27054 21094 27254
rect 21094 27054 21109 27254
rect 22109 27230 22118 27530
rect 22118 27230 22152 27530
rect 22152 27230 22161 27530
rect 23161 27330 23176 27530
rect 23176 27330 23210 27530
rect 23210 27330 23225 27530
rect 24225 27230 24234 27530
rect 24234 27230 24268 27530
rect 24268 27230 24277 27530
rect 21450 26995 22090 27004
rect 21450 26961 22090 26995
rect 21450 26952 22090 26961
rect 22508 26995 23148 27004
rect 23566 26995 24206 27005
rect 25277 27054 25292 27254
rect 25292 27054 25326 27254
rect 25326 27054 25341 27254
rect 22508 26961 23148 26995
rect 23566 26961 24206 26995
rect 22508 26952 23148 26961
rect 23566 26953 24206 26961
rect 24624 26995 25264 27004
rect 24624 26961 25264 26995
rect 24624 26952 25264 26961
rect 25546 26979 25643 27793
rect 21990 26756 22090 26856
rect 22180 26756 22280 26856
rect 23238 26756 23338 26856
rect 25164 26756 25264 26856
rect 21122 26574 21222 26674
rect 23048 26574 23148 26674
rect 24106 26574 24206 26674
rect 24296 26574 24396 26674
rect 21122 26461 21762 26470
rect 21122 26427 21762 26461
rect 21122 26418 21762 26427
rect 22180 26461 22820 26470
rect 23238 26461 23878 26470
rect 22180 26427 22820 26461
rect 23238 26427 23878 26461
rect 22180 26418 22820 26427
rect 21045 26168 21060 26368
rect 21060 26168 21094 26368
rect 21094 26168 21109 26368
rect 22109 25892 22118 26192
rect 22118 25892 22152 26192
rect 22152 25892 22161 26192
rect 23238 26418 23878 26427
rect 24296 26461 24936 26470
rect 24296 26427 24936 26461
rect 24296 26418 24936 26427
rect 23161 25892 23176 26092
rect 23176 25892 23210 26092
rect 23210 25892 23225 26092
rect 24225 25892 24234 26192
rect 24234 25892 24268 26192
rect 24268 25892 24277 26192
rect 25277 26168 25292 26368
rect 25292 26168 25326 26368
rect 25326 26168 25341 26368
rect 20762 25500 25311 25590
rect 20797 25493 25311 25500
rect 16685 25215 18748 25451
rect 11872 24884 12019 24892
rect 11872 24883 12148 24884
rect 19692 24883 19698 24929
rect 19698 24883 19814 24929
rect 11872 24780 19814 24883
rect 11872 23590 12019 24780
rect 19692 24768 19698 24780
rect 19698 24768 19814 24780
rect 19814 24768 19839 24929
rect 19692 24746 19839 24768
rect 22120 25257 24248 25360
rect 22120 24719 22178 25257
rect 12133 24413 12148 24513
rect 12148 24413 12182 24513
rect 12182 24413 12197 24513
rect 14077 24413 14086 24513
rect 14086 24413 14120 24513
rect 14120 24413 14129 24513
rect 16009 24237 16024 24337
rect 16024 24237 16058 24337
rect 16058 24237 16073 24337
rect 17953 24413 17962 24513
rect 17962 24413 17996 24513
rect 17996 24413 18005 24513
rect 22213 24517 22245 24654
rect 22245 24517 22279 24654
rect 22279 24517 22307 24654
rect 19885 24413 19900 24513
rect 19900 24413 19934 24513
rect 19934 24413 19949 24513
rect 22694 24923 22703 25083
rect 22703 24923 22737 25083
rect 22737 24923 22746 25083
rect 23132 24775 23161 24912
rect 23161 24775 23195 24912
rect 23195 24775 23226 24912
rect 23610 24923 23619 25083
rect 23619 24923 23653 25083
rect 23653 24923 23662 25083
rect 24048 24517 24077 24654
rect 24077 24517 24111 24654
rect 24111 24517 24142 24654
rect 22475 24457 22675 24466
rect 22475 24423 22675 24457
rect 22475 24414 22675 24423
rect 22933 24457 23133 24466
rect 22933 24423 23133 24457
rect 22933 24414 23133 24423
rect 23391 24457 23591 24466
rect 23391 24423 23591 24457
rect 23391 24414 23591 24423
rect 23849 24457 24049 24466
rect 23849 24423 24049 24457
rect 23849 24414 24049 24423
rect 20736 24242 20819 24342
rect 22575 24242 22675 24342
rect 22765 24242 22865 24342
rect 23223 24242 23323 24342
rect 23949 24242 24049 24342
rect 12133 23827 12148 23927
rect 12148 23827 12182 23927
rect 12182 23827 12197 23927
rect 14077 23827 14086 23927
rect 14086 23827 14120 23927
rect 14120 23827 14129 23927
rect 16009 24003 16024 24103
rect 16024 24003 16058 24103
rect 16058 24003 16073 24103
rect 17953 23827 17962 23927
rect 17962 23827 17996 23927
rect 17996 23827 18005 23927
rect 20726 24056 20839 24156
rect 22307 24056 22407 24156
rect 23033 24056 23133 24156
rect 23491 24056 23591 24156
rect 23681 24056 23781 24156
rect 19885 23827 19900 23927
rect 19900 23827 19934 23927
rect 19934 23827 19949 23927
rect 22307 23960 22507 23969
rect 22307 23926 22507 23960
rect 22307 23917 22507 23926
rect 22765 23960 22965 23969
rect 22765 23926 22965 23960
rect 22765 23917 22965 23926
rect 23223 23960 23423 23969
rect 23223 23926 23423 23960
rect 23223 23917 23423 23926
rect 23681 23960 23881 23969
rect 23681 23926 23881 23960
rect 23681 23917 23881 23926
rect 22214 23728 22245 23865
rect 22245 23728 22279 23865
rect 22279 23728 22308 23865
rect 11872 23589 12113 23590
rect 11872 23392 19791 23589
rect 22111 23052 22185 23683
rect 22694 23300 22703 23460
rect 22703 23300 22737 23460
rect 22737 23300 22746 23460
rect 23131 23517 23161 23654
rect 23161 23517 23195 23654
rect 23195 23517 23225 23654
rect 23610 23300 23619 23460
rect 23619 23300 23653 23460
rect 23653 23300 23662 23460
rect 24046 23728 24077 23865
rect 24077 23728 24111 23865
rect 24111 23728 24140 23865
rect 25207 24334 25311 25493
rect 25384 24765 25393 24965
rect 25393 24765 25427 24965
rect 25427 24765 25436 24965
rect 25740 24765 25749 24965
rect 25749 24765 25783 24965
rect 25783 24765 25792 24965
rect 25512 24469 25521 24669
rect 25521 24469 25555 24669
rect 25555 24469 25564 24669
rect 25868 24469 25877 24669
rect 25877 24469 25911 24669
rect 25911 24469 25920 24669
rect 25512 24004 25564 24083
rect 25424 23784 25433 23855
rect 25433 23784 25467 23855
rect 25467 23784 25476 23855
rect 25868 23889 25877 23960
rect 25877 23889 25911 23960
rect 25911 23889 25920 23960
rect 25780 23784 25789 23855
rect 25789 23784 25823 23855
rect 25823 23784 25832 23855
rect 24611 23228 25989 23500
rect 17324 22485 17475 22497
rect 12053 15122 12227 21700
rect 12478 21570 12678 21585
rect 12478 21536 12678 21570
rect 14535 21570 14735 21579
rect 12478 21521 12678 21536
rect 13295 21408 13304 21508
rect 13304 21408 13338 21508
rect 13338 21408 13347 21508
rect 13521 21456 13573 21556
rect 13054 21312 13254 21323
rect 13054 21278 13254 21312
rect 13054 21267 13254 21278
rect 13521 21198 13573 21298
rect 12830 21054 12930 21063
rect 12830 21020 12930 21054
rect 12830 21011 12930 21020
rect 12824 20882 12929 20934
rect 13295 20892 13304 20992
rect 13304 20892 13338 20992
rect 13338 20892 13347 20992
rect 12478 20796 12678 20805
rect 12478 20762 12678 20796
rect 12478 20753 12678 20762
rect 12827 20620 12927 20672
rect 12830 20538 12930 20547
rect 12830 20504 12930 20538
rect 12830 20495 12930 20504
rect 13295 20351 13304 20476
rect 13304 20351 13338 20476
rect 13338 20351 13347 20476
rect 13521 20424 13573 20524
rect 13054 20280 13254 20291
rect 13054 20246 13254 20280
rect 13054 20235 13254 20246
rect 12478 20022 12678 20037
rect 12478 19988 12678 20022
rect 12478 19973 12678 19988
rect 13054 19764 13254 19775
rect 13054 19730 13254 19764
rect 13054 19719 13254 19730
rect 13521 19650 13573 19750
rect 12830 19506 12930 19515
rect 12830 19472 12930 19506
rect 12830 19463 12930 19472
rect 12829 19329 12929 19381
rect 13295 19344 13304 19444
rect 13304 19344 13338 19444
rect 13338 19344 13347 19444
rect 12478 19248 12678 19256
rect 12478 19214 12678 19248
rect 12478 19204 12678 19214
rect 12832 19077 12932 19129
rect 12830 18990 12930 18999
rect 12830 18956 12930 18990
rect 12830 18947 12930 18956
rect 13295 18802 13304 18928
rect 13304 18802 13338 18928
rect 13338 18802 13347 18928
rect 13521 18876 13573 18976
rect 13054 18732 13254 18743
rect 13054 18698 13254 18732
rect 13054 18687 13254 18698
rect 12478 18474 12678 18489
rect 12478 18440 12678 18474
rect 12478 18425 12678 18440
rect 13054 18216 13254 18227
rect 13054 18182 13254 18216
rect 13054 18171 13254 18182
rect 13521 18102 13573 18202
rect 12830 17958 12930 17967
rect 12830 17924 12930 17958
rect 12830 17915 12930 17924
rect 12831 17784 12931 17836
rect 13295 17796 13304 17896
rect 13304 17796 13338 17896
rect 13338 17796 13347 17896
rect 12478 17700 12678 17709
rect 12478 17666 12678 17700
rect 12478 17657 12678 17666
rect 12829 17522 12929 17574
rect 12830 17442 12930 17451
rect 12830 17408 12930 17442
rect 12830 17399 12930 17408
rect 13295 17254 13304 17380
rect 13304 17254 13338 17380
rect 13338 17254 13347 17380
rect 13521 17328 13573 17428
rect 13054 17184 13254 17195
rect 13054 17150 13254 17184
rect 13054 17139 13254 17150
rect 12478 16926 12678 16941
rect 12478 16892 12678 16926
rect 12478 16877 12678 16892
rect 13054 16668 13254 16679
rect 13054 16634 13254 16668
rect 13054 16623 13254 16634
rect 13521 16554 13573 16654
rect 12830 16410 12930 16419
rect 12830 16376 12930 16410
rect 12830 16367 12930 16376
rect 12830 16240 12930 16292
rect 13295 16248 13304 16348
rect 13304 16248 13338 16348
rect 13338 16248 13347 16348
rect 12478 16152 12678 16161
rect 12478 16118 12678 16152
rect 12478 16109 12678 16118
rect 12830 15975 12930 16027
rect 12830 15894 12930 15903
rect 12830 15860 12930 15894
rect 12830 15851 12930 15860
rect 13295 15732 13304 15832
rect 13304 15732 13338 15832
rect 13338 15732 13347 15832
rect 13521 15780 13573 15880
rect 13054 15636 13254 15647
rect 13054 15602 13254 15636
rect 13054 15591 13254 15602
rect 12478 15378 12678 15393
rect 12478 15344 12678 15378
rect 12478 15329 12678 15344
rect 13666 21456 13718 21556
rect 14535 21536 14735 21570
rect 14535 21527 14735 21536
rect 13866 21408 13875 21508
rect 13875 21408 13909 21508
rect 13909 21408 13918 21508
rect 14258 21395 14358 21447
rect 14260 21312 14360 21321
rect 14260 21278 14360 21312
rect 14260 21269 14360 21278
rect 13866 21082 13875 21250
rect 13875 21082 13909 21250
rect 13909 21082 13918 21250
rect 13866 21066 13918 21082
rect 13666 20940 13718 21040
rect 14535 21054 14735 21065
rect 14535 21020 14735 21054
rect 14535 21009 14735 21020
rect 13959 20796 14159 20811
rect 13959 20762 14159 20796
rect 13959 20747 14159 20762
rect 14535 20538 14735 20549
rect 14535 20504 14735 20538
rect 14535 20493 14735 20504
rect 13666 20166 13718 20266
rect 14260 20280 14360 20289
rect 14260 20246 14360 20280
rect 14260 20237 14360 20246
rect 13866 20118 13875 20218
rect 13875 20118 13909 20218
rect 13909 20118 13918 20218
rect 14260 20103 14360 20155
rect 14535 20022 14735 20031
rect 14535 19988 14735 20022
rect 14535 19979 14735 19988
rect 14262 19848 14362 19900
rect 14260 19764 14360 19773
rect 14260 19730 14360 19764
rect 14260 19721 14360 19730
rect 13866 19534 13875 19702
rect 13875 19534 13909 19702
rect 13909 19534 13918 19702
rect 13866 19518 13918 19534
rect 13666 19392 13718 19492
rect 14535 19506 14735 19517
rect 14535 19472 14735 19506
rect 14535 19461 14735 19472
rect 13959 19248 14159 19263
rect 13959 19214 14159 19248
rect 13959 19199 14159 19214
rect 14535 18990 14735 19001
rect 14535 18956 14735 18990
rect 14535 18945 14735 18956
rect 13666 18618 13718 18718
rect 14259 18732 14359 18741
rect 14259 18698 14359 18732
rect 14259 18689 14359 18698
rect 13866 18570 13875 18670
rect 13875 18570 13909 18670
rect 13909 18570 13918 18670
rect 14262 18552 14362 18604
rect 14535 18474 14735 18483
rect 14535 18440 14735 18474
rect 14535 18431 14735 18440
rect 14260 18290 14360 18342
rect 14260 18216 14360 18225
rect 14260 18182 14360 18216
rect 14260 18173 14360 18182
rect 13866 17986 13875 18154
rect 13875 17986 13909 18154
rect 13909 17986 13918 18154
rect 13866 17970 13918 17986
rect 13666 17844 13718 17944
rect 14535 17958 14735 17969
rect 14535 17924 14735 17958
rect 14535 17913 14735 17924
rect 13959 17700 14159 17715
rect 13959 17666 14159 17700
rect 13959 17651 14159 17666
rect 14535 17442 14735 17453
rect 14535 17408 14735 17442
rect 14535 17397 14735 17408
rect 13666 17070 13718 17170
rect 14260 17184 14360 17193
rect 14260 17150 14360 17184
rect 14260 17141 14360 17150
rect 13866 17022 13875 17122
rect 13875 17022 13909 17122
rect 13909 17022 13918 17122
rect 14258 17004 14358 17056
rect 14535 16926 14735 16935
rect 14535 16892 14735 16926
rect 14535 16883 14735 16892
rect 14259 16748 14359 16800
rect 14260 16668 14360 16677
rect 14260 16634 14360 16668
rect 14260 16625 14360 16634
rect 13866 16438 13875 16606
rect 13875 16438 13909 16606
rect 13909 16438 13918 16606
rect 13866 16406 13918 16438
rect 14535 16410 14735 16421
rect 13666 16296 13718 16396
rect 14535 16376 14735 16410
rect 14535 16365 14735 16376
rect 13959 16152 14159 16167
rect 13959 16118 14159 16152
rect 13959 16103 14159 16118
rect 14534 15894 14734 15905
rect 14534 15860 14734 15894
rect 14534 15849 14734 15860
rect 13666 15522 13718 15622
rect 14260 15636 14360 15645
rect 14260 15602 14360 15636
rect 14260 15593 14360 15602
rect 13866 15474 13875 15574
rect 13875 15474 13909 15574
rect 13909 15474 13918 15574
rect 14262 15470 14362 15522
rect 14535 15378 14735 15387
rect 14535 15344 14735 15378
rect 14535 15335 14735 15344
rect 14994 15315 15106 21656
rect 15736 17060 15927 22467
rect 16883 22440 17006 22449
rect 16883 22406 17006 22440
rect 16883 22397 17006 22406
rect 16096 22375 16156 22384
rect 16212 22375 16272 22384
rect 16096 22341 16156 22375
rect 16212 22341 16272 22375
rect 16096 22332 16156 22341
rect 16212 22332 16272 22341
rect 16212 22117 16272 22126
rect 16212 22083 16272 22117
rect 16212 22074 16272 22083
rect 16096 21859 16156 21868
rect 16096 21825 16156 21859
rect 16096 21816 16156 21825
rect 16212 21601 16272 21610
rect 16212 21567 16272 21601
rect 16212 21558 16272 21567
rect 16096 21343 16156 21352
rect 16096 21309 16156 21343
rect 16096 21300 16156 21309
rect 16936 21982 17059 21991
rect 16936 21948 17059 21982
rect 16936 21939 17059 21948
rect 16883 21859 17006 21868
rect 16883 21825 17006 21859
rect 16883 21816 17006 21825
rect 16096 21085 16156 21094
rect 16096 21051 16156 21085
rect 16096 21042 16156 21051
rect 16212 20827 16272 20836
rect 16212 20793 16272 20827
rect 16212 20784 16272 20793
rect 16096 20569 16156 20578
rect 16096 20535 16156 20569
rect 16096 20526 16156 20535
rect 16212 20311 16272 20320
rect 16212 20277 16272 20311
rect 16212 20268 16272 20277
rect 16096 20053 16156 20062
rect 16096 20019 16156 20053
rect 16096 20010 16156 20019
rect 16935 21401 17059 21410
rect 16935 21367 17059 21401
rect 16935 21358 17059 21367
rect 17324 21143 17330 22485
rect 16883 20569 16996 20578
rect 16883 20535 16996 20569
rect 16883 20526 16996 20535
rect 16096 19795 16156 19804
rect 16096 19761 16156 19795
rect 16096 19752 16156 19761
rect 16212 19537 16272 19546
rect 16212 19503 16272 19537
rect 16212 19494 16272 19503
rect 16096 19279 16156 19288
rect 16096 19245 16156 19279
rect 16096 19236 16156 19245
rect 16212 19021 16272 19030
rect 16212 18987 16272 19021
rect 16212 18978 16272 18987
rect 16096 18763 16156 18772
rect 16096 18729 16156 18763
rect 16096 18720 16156 18729
rect 16936 20111 17059 20120
rect 16936 20077 17059 20111
rect 16936 20068 17059 20077
rect 16883 19279 16996 19288
rect 16883 19245 16996 19279
rect 16883 19236 16996 19245
rect 16096 18505 16156 18514
rect 16096 18471 16156 18505
rect 16096 18462 16156 18471
rect 16212 18247 16272 18256
rect 16212 18213 16272 18247
rect 16212 18204 16272 18213
rect 16096 17989 16156 17998
rect 16096 17955 16156 17989
rect 16096 17946 16156 17955
rect 16212 17731 16272 17740
rect 16212 17697 16272 17731
rect 16212 17688 16272 17697
rect 16096 17473 16156 17482
rect 16096 17439 16156 17473
rect 16096 17430 16156 17439
rect 16936 18821 17059 18830
rect 16936 18787 17059 18821
rect 16936 18778 17059 18787
rect 16883 17989 16996 17998
rect 16883 17955 16996 17989
rect 16883 17946 16996 17955
rect 16096 17215 16156 17224
rect 16096 17181 16156 17215
rect 16096 17172 16156 17181
rect 16936 17531 17059 17540
rect 16936 17497 17059 17531
rect 16936 17488 17059 17497
rect 17330 17490 17469 22485
rect 17469 21143 17475 22485
rect 22066 23045 22293 23052
rect 22066 22882 23409 23045
rect 22066 21866 22404 22882
rect 22404 22875 23409 22882
rect 23333 22750 23742 22766
rect 23333 22716 23742 22750
rect 23333 22701 23742 22716
rect 22571 22533 22582 22673
rect 22582 22533 22616 22673
rect 22616 22533 22627 22673
rect 22666 22392 23166 22407
rect 22666 22358 23166 22392
rect 22666 22343 23166 22358
rect 23333 22034 23742 22050
rect 23333 22000 23742 22034
rect 23333 21985 23742 22000
rect 23955 21866 24166 22917
rect 24907 23000 25109 23008
rect 24907 22962 25109 23000
rect 24907 22956 25109 22962
rect 25741 23000 25943 23007
rect 25741 22962 25943 23000
rect 25741 22955 25943 22962
rect 22066 21627 24166 21866
rect 22066 21625 22293 21627
rect 23955 21616 24166 21627
rect 16883 16901 17023 16916
rect 16883 16867 17023 16901
rect 16883 16852 17023 16867
rect 16919 16643 17059 16652
rect 16919 16609 17059 16643
rect 16919 16600 17059 16609
rect 15334 16208 16377 16316
rect 16883 16385 17023 16400
rect 16883 16351 17023 16385
rect 16883 16336 17023 16351
rect 15580 16008 16180 16015
rect 15580 15974 15620 16008
rect 15620 15974 15654 16008
rect 15654 15974 15720 16008
rect 15720 15974 15754 16008
rect 15754 15974 15820 16008
rect 15820 15974 15854 16008
rect 15854 15974 15920 16008
rect 15920 15974 15954 16008
rect 15954 15974 16020 16008
rect 16020 15974 16054 16008
rect 16054 15974 16120 16008
rect 16120 15974 16154 16008
rect 16154 15974 16180 16008
rect 15580 15941 16180 15974
rect 15155 15307 15251 15834
rect 12309 15125 12461 15179
rect 13299 15125 13447 15179
rect 15767 15161 16246 15281
rect 16344 15258 16492 16083
rect 16763 15749 16790 16108
rect 16790 15749 16824 16108
rect 16824 15749 16828 16108
rect 17216 16941 17251 17028
rect 17251 16941 17351 17028
rect 17216 16042 17351 16941
rect 16883 15718 16959 15727
rect 16883 15684 16959 15718
rect 16883 15675 16959 15684
rect 16763 15295 16790 15654
rect 16790 15295 16824 15654
rect 16824 15295 16828 15654
rect 17218 15049 17350 16042
rect 17429 15050 17577 17029
rect 17910 11015 25708 11104
rect 2688 3829 2862 10407
rect 2944 10350 3096 10404
rect 3934 10350 4082 10404
rect 3113 10185 3313 10200
rect 3113 10151 3313 10185
rect 3113 10136 3313 10151
rect 3689 9927 3889 9938
rect 3689 9893 3889 9927
rect 3689 9882 3889 9893
rect 3930 9697 3939 9797
rect 3939 9697 3973 9797
rect 3973 9697 3982 9797
rect 5170 10185 5370 10194
rect 5170 10151 5370 10185
rect 5170 10142 5370 10151
rect 3465 9669 3565 9678
rect 3465 9635 3565 9669
rect 3465 9626 3565 9635
rect 4156 9649 4208 9749
rect 3465 9502 3565 9554
rect 3113 9411 3313 9420
rect 3113 9377 3313 9411
rect 3113 9368 3313 9377
rect 3465 9237 3565 9289
rect 3930 9181 3939 9281
rect 3939 9181 3973 9281
rect 3973 9181 3982 9281
rect 3465 9153 3565 9162
rect 3465 9119 3565 9153
rect 3465 9110 3565 9119
rect 3689 8895 3889 8906
rect 3689 8861 3889 8895
rect 3689 8850 3889 8861
rect 3113 8637 3313 8652
rect 3113 8603 3313 8637
rect 3113 8588 3313 8603
rect 3689 8379 3889 8390
rect 3689 8345 3889 8379
rect 3689 8334 3889 8345
rect 4156 8875 4208 8975
rect 3930 8149 3939 8275
rect 3939 8149 3973 8275
rect 3973 8149 3982 8275
rect 3465 8121 3565 8130
rect 3465 8087 3565 8121
rect 3465 8078 3565 8087
rect 4156 8101 4208 8201
rect 3464 7955 3564 8007
rect 3113 7863 3313 7872
rect 3113 7829 3313 7863
rect 3113 7820 3313 7829
rect 3466 7693 3566 7745
rect 3930 7633 3939 7733
rect 3939 7633 3973 7733
rect 3973 7633 3982 7733
rect 3465 7605 3565 7614
rect 3465 7571 3565 7605
rect 3465 7562 3565 7571
rect 3689 7347 3889 7358
rect 3689 7313 3889 7347
rect 3689 7302 3889 7313
rect 3113 7089 3313 7104
rect 3113 7055 3313 7089
rect 3113 7040 3313 7055
rect 3689 6831 3889 6842
rect 3689 6797 3889 6831
rect 3689 6786 3889 6797
rect 4156 7327 4208 7427
rect 3930 6601 3939 6727
rect 3939 6601 3973 6727
rect 3973 6601 3982 6727
rect 3465 6573 3565 6582
rect 3465 6539 3565 6573
rect 3465 6530 3565 6539
rect 4156 6553 4208 6653
rect 3467 6400 3567 6452
rect 3113 6315 3313 6325
rect 3113 6281 3313 6315
rect 3113 6273 3313 6281
rect 3464 6148 3564 6200
rect 3930 6085 3939 6185
rect 3939 6085 3973 6185
rect 3973 6085 3982 6185
rect 3465 6057 3565 6066
rect 3465 6023 3565 6057
rect 3465 6014 3565 6023
rect 3689 5799 3889 5810
rect 3689 5765 3889 5799
rect 3689 5754 3889 5765
rect 3113 5541 3313 5556
rect 3113 5507 3313 5541
rect 3113 5492 3313 5507
rect 3689 5283 3889 5294
rect 3689 5249 3889 5283
rect 3689 5238 3889 5249
rect 4156 5779 4208 5879
rect 3930 5053 3939 5178
rect 3939 5053 3973 5178
rect 3973 5053 3982 5178
rect 3465 5025 3565 5034
rect 3465 4991 3565 5025
rect 3465 4982 3565 4991
rect 4156 5005 4208 5105
rect 3462 4857 3562 4909
rect 3113 4767 3313 4776
rect 3113 4733 3313 4767
rect 3113 4724 3313 4733
rect 3459 4595 3564 4647
rect 3930 4537 3939 4637
rect 3939 4537 3973 4637
rect 3973 4537 3982 4637
rect 3465 4509 3565 4518
rect 3465 4475 3565 4509
rect 3465 4466 3565 4475
rect 3689 4251 3889 4262
rect 3689 4217 3889 4251
rect 3689 4206 3889 4217
rect 4156 4231 4208 4331
rect 3930 4021 3939 4121
rect 3939 4021 3973 4121
rect 3973 4021 3982 4121
rect 3113 3993 3313 4008
rect 3113 3959 3313 3993
rect 4156 3973 4208 4073
rect 4301 9907 4353 10007
rect 4501 9955 4510 10055
rect 4510 9955 4544 10055
rect 4544 9955 4553 10055
rect 4897 10007 4997 10059
rect 4895 9927 4995 9936
rect 4895 9893 4995 9927
rect 4895 9884 4995 9893
rect 4301 9133 4353 9233
rect 5169 9669 5369 9680
rect 5169 9635 5369 9669
rect 5169 9624 5369 9635
rect 4594 9411 4794 9426
rect 4594 9377 4794 9411
rect 4594 9362 4794 9377
rect 5170 9153 5370 9164
rect 4501 9091 4553 9123
rect 5170 9119 5370 9153
rect 5170 9108 5370 9119
rect 4501 8923 4510 9091
rect 4510 8923 4544 9091
rect 4544 8923 4553 9091
rect 4895 8895 4995 8904
rect 4895 8861 4995 8895
rect 4895 8852 4995 8861
rect 4894 8729 4994 8781
rect 5170 8637 5370 8646
rect 5170 8603 5370 8637
rect 5170 8594 5370 8603
rect 4301 8359 4353 8459
rect 4501 8407 4510 8507
rect 4510 8407 4544 8507
rect 4544 8407 4553 8507
rect 4893 8473 4993 8525
rect 4895 8379 4995 8388
rect 4895 8345 4995 8379
rect 4895 8336 4995 8345
rect 4301 7585 4353 7685
rect 5170 8121 5370 8132
rect 5170 8087 5370 8121
rect 5170 8076 5370 8087
rect 4594 7863 4794 7878
rect 4594 7829 4794 7863
rect 4594 7814 4794 7829
rect 5170 7605 5370 7616
rect 5170 7571 5370 7605
rect 4501 7543 4553 7559
rect 5170 7560 5370 7571
rect 4501 7375 4510 7543
rect 4510 7375 4544 7543
rect 4544 7375 4553 7543
rect 4895 7347 4995 7356
rect 4895 7313 4995 7347
rect 4895 7304 4995 7313
rect 4895 7187 4995 7239
rect 5170 7089 5370 7098
rect 5170 7055 5370 7089
rect 5170 7046 5370 7055
rect 4301 6811 4353 6911
rect 4501 6859 4510 6959
rect 4510 6859 4544 6959
rect 4544 6859 4553 6959
rect 4897 6925 4997 6977
rect 4894 6831 4994 6840
rect 4894 6797 4994 6831
rect 4894 6788 4994 6797
rect 4301 6037 4353 6137
rect 5170 6573 5370 6584
rect 5170 6539 5370 6573
rect 5170 6528 5370 6539
rect 4594 6315 4794 6330
rect 4594 6281 4794 6315
rect 4594 6266 4794 6281
rect 5170 6057 5370 6068
rect 5170 6023 5370 6057
rect 4501 5995 4553 6011
rect 5170 6012 5370 6023
rect 4501 5827 4510 5995
rect 4510 5827 4544 5995
rect 4544 5827 4553 5995
rect 4895 5799 4995 5808
rect 4895 5765 4995 5799
rect 4895 5756 4995 5765
rect 4897 5629 4997 5681
rect 5170 5541 5370 5550
rect 5170 5507 5370 5541
rect 5170 5498 5370 5507
rect 4301 5263 4353 5363
rect 4501 5311 4510 5411
rect 4510 5311 4544 5411
rect 4544 5311 4553 5411
rect 4895 5374 4995 5426
rect 4895 5283 4995 5292
rect 4895 5249 4995 5283
rect 4895 5240 4995 5249
rect 4301 4489 4353 4589
rect 5170 5025 5370 5036
rect 5170 4991 5370 5025
rect 5170 4980 5370 4991
rect 4594 4767 4794 4782
rect 4594 4733 4794 4767
rect 4594 4718 4794 4733
rect 5170 4509 5370 4520
rect 5170 4475 5370 4509
rect 4501 4447 4553 4463
rect 5170 4464 5370 4475
rect 4501 4279 4510 4447
rect 4510 4279 4544 4447
rect 4544 4279 4553 4447
rect 4895 4251 4995 4260
rect 4895 4217 4995 4251
rect 4895 4208 4995 4217
rect 4301 3973 4353 4073
rect 4501 4021 4510 4121
rect 4510 4021 4544 4121
rect 4544 4021 4553 4121
rect 4893 4082 4993 4134
rect 5170 3993 5370 4002
rect 3113 3944 3313 3959
rect 5170 3959 5370 3993
rect 5170 3950 5370 3959
rect 5629 3873 5741 10214
rect 5790 9695 5886 10222
rect 6402 10248 6881 10368
rect 6215 9555 6815 9588
rect 6215 9521 6255 9555
rect 6255 9521 6289 9555
rect 6289 9521 6355 9555
rect 6355 9521 6389 9555
rect 6389 9521 6455 9555
rect 6455 9521 6489 9555
rect 6489 9521 6555 9555
rect 6555 9521 6589 9555
rect 6589 9521 6655 9555
rect 6655 9521 6689 9555
rect 6689 9521 6755 9555
rect 6755 9521 6789 9555
rect 6789 9521 6815 9555
rect 6215 9514 6815 9521
rect 6979 9446 7127 10271
rect 7398 9875 7425 10234
rect 7425 9875 7459 10234
rect 7459 9875 7463 10234
rect 7518 9845 7594 9854
rect 7518 9811 7594 9845
rect 7518 9802 7594 9811
rect 7398 9421 7425 9780
rect 7425 9421 7459 9780
rect 7459 9421 7463 9780
rect 7853 9487 7985 10480
rect 5969 9213 7012 9321
rect 7518 9178 7658 9193
rect 7518 9144 7658 9178
rect 7518 9129 7658 9144
rect 7554 8920 7694 8929
rect 7554 8886 7694 8920
rect 7554 8877 7694 8886
rect 6371 2963 6562 8370
rect 6731 8249 6791 8258
rect 6731 8215 6791 8249
rect 6731 8206 6791 8215
rect 6731 7991 6791 8000
rect 6731 7957 6791 7991
rect 6731 7948 6791 7957
rect 6847 7733 6907 7742
rect 6847 7699 6907 7733
rect 6847 7690 6907 7699
rect 6731 7475 6791 7484
rect 6731 7441 6791 7475
rect 6731 7432 6791 7441
rect 6847 7217 6907 7226
rect 6847 7183 6907 7217
rect 6847 7174 6907 7183
rect 7518 8662 7658 8677
rect 7518 8628 7658 8662
rect 7518 8613 7658 8628
rect 7851 8588 7986 9487
rect 7851 8501 7886 8588
rect 7886 8501 7986 8588
rect 8064 8500 8212 10479
rect 21823 10318 21833 10654
rect 21833 10318 21867 10654
rect 21867 10318 21877 10654
rect 18142 9830 18175 10135
rect 18175 9830 18209 10135
rect 18209 9830 18218 10135
rect 21823 9830 21833 10166
rect 21833 9830 21867 10166
rect 21867 9830 21877 10166
rect 25483 9830 25491 10125
rect 25491 9830 25525 10125
rect 25525 9830 25559 10125
rect 18142 9368 18451 9452
rect 18950 9377 19299 9444
rect 24014 9374 24363 9441
rect 26498 9298 26678 9459
rect 19377 9187 19726 9254
rect 24434 9191 24783 9258
rect 25148 9188 25538 9258
rect 19341 8214 19385 8782
rect 19385 8214 19419 8782
rect 19419 8214 19427 8782
rect 7571 7933 7694 7942
rect 7571 7899 7694 7933
rect 7571 7890 7694 7899
rect 6731 6959 6791 6968
rect 6731 6925 6791 6959
rect 6731 6916 6791 6925
rect 6731 6701 6791 6710
rect 6731 6667 6791 6701
rect 6731 6658 6791 6667
rect 6847 6443 6907 6452
rect 6847 6409 6907 6443
rect 6847 6400 6907 6409
rect 6731 6185 6791 6194
rect 6731 6151 6791 6185
rect 6731 6142 6791 6151
rect 6847 5927 6907 5936
rect 6847 5893 6907 5927
rect 6847 5884 6907 5893
rect 7518 7475 7631 7484
rect 7518 7441 7631 7475
rect 7518 7432 7631 7441
rect 7571 6643 7694 6652
rect 7571 6609 7694 6643
rect 7571 6600 7694 6609
rect 6731 5669 6791 5678
rect 6731 5635 6791 5669
rect 6731 5626 6791 5635
rect 6731 5411 6791 5420
rect 6731 5377 6791 5411
rect 6731 5368 6791 5377
rect 6847 5153 6907 5162
rect 6847 5119 6907 5153
rect 6847 5110 6907 5119
rect 6731 4895 6791 4904
rect 6731 4861 6791 4895
rect 6731 4852 6791 4861
rect 6847 4637 6907 4646
rect 6847 4603 6907 4637
rect 6847 4594 6907 4603
rect 7518 6185 7631 6194
rect 7518 6151 7631 6185
rect 7518 6142 7631 6151
rect 7571 5353 7694 5362
rect 7571 5319 7694 5353
rect 7571 5310 7694 5319
rect 6731 4379 6791 4388
rect 6731 4345 6791 4379
rect 6731 4336 6791 4345
rect 6731 4121 6791 4130
rect 6731 4087 6791 4121
rect 6731 4078 6791 4087
rect 6847 3863 6907 3872
rect 6847 3829 6907 3863
rect 6847 3820 6907 3829
rect 6731 3605 6791 3614
rect 6731 3571 6791 3605
rect 6731 3562 6791 3571
rect 6847 3347 6907 3356
rect 6847 3313 6907 3347
rect 6847 3304 6907 3313
rect 6731 3089 6791 3098
rect 7518 4895 7631 4904
rect 7518 4861 7631 4895
rect 7518 4852 7631 4861
rect 7570 4063 7694 4072
rect 7570 4029 7694 4063
rect 7570 4020 7694 4029
rect 7518 3605 7641 3614
rect 7518 3571 7641 3605
rect 7518 3562 7641 3571
rect 7571 3482 7694 3491
rect 7571 3448 7694 3482
rect 7571 3439 7694 3448
rect 6847 3089 6907 3098
rect 6731 3055 6791 3089
rect 6847 3055 6907 3089
rect 6731 3046 6791 3055
rect 6847 3046 6907 3055
rect 7518 3024 7641 3033
rect 7518 2990 7641 3024
rect 7518 2981 7641 2990
rect 7959 2945 7965 4287
rect 7965 2945 8104 7940
rect 21835 7638 21843 7957
rect 21843 7638 21877 7957
rect 21877 7638 21887 7957
rect 24293 8214 24301 8782
rect 24301 8214 24335 8782
rect 24335 8214 24379 8782
rect 19451 7556 19661 7568
rect 19451 7522 19661 7556
rect 19451 7511 19661 7522
rect 24063 7556 24273 7568
rect 24063 7522 24273 7556
rect 24063 7511 24273 7522
rect 19474 7393 19661 7450
rect 21904 7390 22105 7454
rect 18058 7269 18634 7286
rect 18058 7235 18634 7269
rect 18058 7231 18634 7235
rect 21604 7078 21814 7135
rect 24063 7080 24273 7137
rect 18676 6239 18684 7038
rect 18684 6239 18718 7038
rect 18718 6239 18728 7038
rect 21604 6991 21814 7003
rect 21604 6957 21814 6991
rect 21604 6946 21814 6957
rect 21904 6991 22114 7002
rect 21904 6957 22114 6991
rect 19274 5835 19384 6907
rect 19384 5835 19418 6907
rect 19418 5835 19426 6907
rect 21904 6945 22114 6957
rect 21834 6557 21842 6876
rect 21842 6557 21876 6876
rect 21876 6557 21886 6876
rect 17832 5573 18385 5667
rect 19446 5681 19926 5688
rect 19446 5647 19926 5681
rect 19446 5636 19926 5647
rect 21904 5681 22384 5689
rect 24291 5835 24300 6907
rect 24300 5835 24334 6907
rect 24334 5835 24443 6907
rect 21904 5647 22384 5681
rect 21904 5637 22384 5647
rect 17834 5343 24768 5432
rect 8104 2945 8110 4287
rect 7959 2933 8110 2945
<< metal2 >>
rect 11711 33012 14392 33022
rect 11711 32798 11800 33012
rect 11712 31193 11800 32798
rect 11238 31191 11800 31193
rect 3217 31121 11800 31191
rect 3217 30961 10935 31121
rect 11665 30961 11800 31121
rect 3217 30890 11800 30961
rect 3217 30801 3401 30890
rect 11199 30801 11800 30890
rect 3217 30791 11800 30801
rect 7314 30440 7368 30791
rect 11238 30790 11800 30791
rect 3623 29921 3709 29964
rect 3623 29616 3633 29921
rect 3623 29248 3709 29616
rect 7314 29952 7368 30104
rect 7314 29606 7368 29616
rect 10974 29911 11060 29964
rect 11050 29616 11060 29911
rect 3623 29238 3942 29248
rect 3623 29154 3633 29238
rect 3623 29144 3942 29154
rect 4441 29230 4802 29245
rect 4790 29163 4802 29230
rect 4441 29145 4802 29163
rect 9505 29227 9870 29245
rect 9854 29160 9870 29227
rect 9505 29145 9870 29160
rect 3549 27082 4125 27092
rect 3549 27007 4125 27017
rect 4167 26833 4219 26834
rect 4164 26824 4222 26833
rect 4164 26823 4167 26824
rect 4219 26823 4222 26824
rect 4164 26015 4222 26025
rect 4716 26703 4802 29145
rect 4832 29040 5218 29060
rect 4832 28973 4868 29040
rect 5217 28973 5218 29040
rect 4832 28960 5218 28973
rect 4832 28568 4918 28960
rect 4832 27990 4918 28000
rect 9784 28568 9870 29145
rect 10974 29060 11060 29616
rect 11965 32799 14392 32809
rect 12557 32516 15238 32526
rect 12629 32426 13433 32516
rect 12557 31906 12629 31916
rect 13505 32426 15238 32516
rect 13433 31906 13505 31916
rect 12999 31777 13063 31787
rect 12999 30767 13063 30777
rect 12122 30540 12186 30550
rect 12122 29530 12186 29540
rect 13875 30540 13939 30550
rect 13875 29530 13939 29540
rect 11800 29391 11965 29401
rect 12200 29490 12480 29500
rect 12200 29428 12480 29438
rect 12638 29490 12918 29500
rect 12638 29428 12918 29438
rect 13076 29490 13356 29500
rect 13076 29428 13356 29438
rect 13514 29490 13794 29500
rect 13514 29428 13794 29438
rect 12200 29245 12300 29428
rect 12200 29135 12300 29145
rect 9784 27990 9870 28000
rect 9900 29044 10274 29060
rect 9900 28977 9925 29044
rect 9900 28960 10274 28977
rect 10639 29044 11060 29060
rect 11029 28974 11060 29044
rect 10639 28960 11060 28974
rect 7322 27756 7378 27766
rect 7322 27404 7378 27414
rect 4942 27354 5152 27364
rect 4942 27236 5152 27297
rect 9554 27354 9764 27364
rect 4942 27179 4965 27236
rect 4942 27169 5152 27179
rect 7395 27240 7605 27252
rect 7596 27176 7605 27240
rect 7095 26921 7305 26931
rect 7095 26789 7305 26864
rect 7095 26722 7305 26732
rect 7395 26788 7605 27176
rect 9554 26923 9764 27297
rect 9554 26856 9764 26866
rect 7395 26721 7605 26731
rect 9900 26703 9986 28960
rect 12448 28936 12548 28946
rect 12448 28651 12548 28836
rect 12638 28936 12738 29428
rect 12638 28826 12738 28836
rect 12886 29245 12986 29255
rect 12886 28651 12986 29145
rect 13076 28936 13176 29428
rect 13076 28826 13176 28836
rect 13324 29245 13424 29255
rect 13324 28651 13424 29145
rect 13514 29245 13614 29428
rect 13514 29135 13614 29145
rect 13762 28936 13862 28946
rect 13762 28651 13862 28836
rect 12268 28641 12548 28651
rect 4716 26693 4917 26703
rect 4716 25621 4765 26693
rect 9782 26693 9986 26703
rect 7321 26672 7379 26682
rect 7321 26323 7379 26333
rect 4917 25621 4919 26129
rect 4716 25552 4919 25621
rect 9934 25621 9986 26693
rect 9782 25611 9986 25621
rect 11817 28583 11965 28593
rect 3015 25519 3113 25529
rect 3113 25453 3997 25519
rect 3113 25359 3323 25453
rect 3876 25359 3997 25453
rect 4937 25477 5417 25487
rect 4937 25409 5417 25419
rect 7395 25479 7875 25489
rect 7395 25411 7875 25421
rect 3113 25228 3997 25359
rect 11816 25407 11817 25417
rect 12268 28579 12548 28589
rect 12706 28641 12986 28651
rect 12706 28579 12986 28589
rect 13144 28641 13424 28651
rect 13144 28579 13424 28589
rect 13582 28641 13862 28651
rect 13582 28579 13862 28589
rect 12123 28539 12187 28549
rect 12123 27529 12187 27539
rect 13875 28539 13939 28549
rect 13875 27529 13939 27539
rect 12999 27379 13063 27389
rect 12999 26369 13063 26379
rect 15138 26995 15238 32426
rect 15329 29245 15621 29255
rect 15329 29135 15621 29145
rect 27028 28171 27326 28181
rect 18739 28167 20751 28171
rect 25689 28169 27028 28170
rect 25642 28168 27028 28169
rect 25403 28167 27028 28168
rect 18739 28158 27028 28167
rect 18739 28157 25403 28158
rect 18739 27792 20700 28157
rect 25662 27793 27028 28158
rect 25504 27792 25546 27793
rect 18739 27781 20762 27792
rect 18739 27508 19138 27781
rect 20692 27753 20762 27781
rect 15475 27498 19138 27508
rect 15475 27197 18851 27207
rect 15138 26985 18682 26995
rect 15138 26895 16958 26985
rect 12557 26173 13957 26174
rect 15138 26173 15238 26895
rect 12557 26163 15238 26173
rect 12629 26074 13432 26163
rect 12557 25553 12629 25563
rect 13504 26074 15238 26163
rect 13829 26073 15238 26074
rect 17010 26895 17794 26985
rect 16958 25975 17010 25985
rect 17376 26609 17428 26619
rect 13432 25553 13504 25563
rect 17846 26895 18630 26985
rect 17794 25975 17846 25985
rect 18212 26609 18264 26619
rect 17376 25461 17428 25609
rect 18630 25975 18682 25985
rect 18851 25681 19138 25691
rect 18212 25461 18264 25609
rect 20879 27783 25546 27792
rect 20879 27782 25504 27783
rect 20879 27753 20907 27782
rect 22109 27530 22161 27782
rect 21045 27254 21109 27264
rect 23161 27530 23225 27540
rect 23161 27320 23225 27330
rect 24225 27530 24277 27782
rect 22109 27220 22161 27230
rect 24225 27220 24277 27230
rect 25277 27254 25341 27264
rect 21045 27044 21109 27054
rect 25277 27044 25341 27054
rect 21450 27004 22090 27014
rect 21450 26942 22090 26952
rect 22508 27004 23148 27014
rect 22508 26942 23148 26952
rect 23566 27005 24206 27015
rect 23566 26943 24206 26953
rect 21990 26856 22090 26942
rect 21990 26746 22090 26756
rect 22180 26856 22280 26866
rect 21122 26674 21222 26684
rect 21122 26480 21222 26574
rect 22180 26480 22280 26756
rect 23048 26674 23148 26942
rect 23048 26564 23148 26574
rect 23238 26856 23338 26866
rect 23238 26480 23338 26756
rect 24106 26674 24206 26943
rect 24624 27004 25264 27014
rect 25643 27784 27028 27793
rect 25643 27783 25662 27784
rect 27028 27774 27326 27784
rect 25546 26969 25643 26979
rect 24624 26942 25264 26952
rect 25164 26856 25264 26942
rect 25164 26746 25264 26756
rect 24106 26564 24206 26574
rect 24296 26674 24396 26684
rect 24296 26480 24396 26574
rect 21122 26470 21762 26480
rect 21122 26408 21762 26418
rect 22180 26470 22820 26480
rect 22180 26408 22820 26418
rect 23238 26470 23878 26480
rect 23238 26408 23878 26418
rect 24296 26470 24936 26480
rect 24296 26408 24936 26418
rect 21045 26368 21109 26378
rect 25277 26368 25341 26378
rect 21045 26158 21109 26168
rect 22109 26192 22161 26202
rect 24225 26192 24277 26202
rect 22109 25600 22161 25892
rect 23161 26092 23225 26102
rect 23161 25882 23225 25892
rect 25277 26158 25341 26168
rect 24225 25600 24277 25892
rect 20879 25590 25311 25600
rect 18838 25565 20450 25575
rect 18962 25506 20450 25565
rect 18838 25496 20450 25506
rect 16685 25451 18748 25461
rect 11965 25374 14381 25384
rect 11816 25230 11929 25231
rect 3113 25218 10259 25228
rect 11816 25221 14381 25230
rect 11929 25220 14381 25221
rect 3113 25129 3325 25218
rect 16685 25205 18748 25215
rect 3113 25119 10259 25129
rect 3015 25109 3113 25119
rect 9850 24895 10259 25119
rect 19692 24929 19839 24939
rect 11872 24895 12019 24902
rect 9847 24894 12019 24895
rect 9847 24893 12148 24894
rect 9847 24892 19692 24893
rect 9847 24558 11872 24892
rect 12019 24884 19692 24892
rect 12148 24883 19692 24884
rect 9129 23600 9383 23610
rect 11870 23600 11872 23604
rect 9383 23594 11872 23600
rect 12019 24770 19692 24780
rect 12133 24513 12197 24523
rect 12133 24403 12197 24413
rect 14077 24513 14129 24770
rect 14077 24403 14129 24413
rect 17953 24513 18005 24770
rect 19692 24736 19839 24746
rect 17953 24403 18005 24413
rect 19885 24513 19949 24523
rect 19885 24403 19949 24413
rect 16009 24337 16073 24347
rect 16009 24227 16073 24237
rect 16009 24103 16073 24113
rect 16009 23993 16073 24003
rect 12133 23927 12197 23937
rect 12133 23817 12197 23827
rect 14077 23927 14129 23937
rect 14077 23604 14129 23827
rect 17953 23927 18005 23937
rect 17953 23604 18005 23827
rect 19885 23927 19949 23937
rect 19885 23817 19949 23827
rect 12019 23599 19325 23604
rect 19859 23599 20043 23609
rect 12019 23594 19859 23599
rect 9383 23391 11870 23594
rect 19325 23589 19859 23594
rect 19791 23392 19859 23589
rect 19325 23391 19859 23392
rect 9383 23382 19859 23391
rect 20043 23382 20052 23599
rect 9129 23372 9383 23382
rect 11870 23381 19325 23382
rect 12042 21700 12237 23381
rect 19859 23372 20043 23382
rect 16576 23071 16676 23081
rect 16576 22678 16676 22891
rect 12042 21514 12053 21700
rect 11526 21341 11683 21351
rect 12043 21341 12053 21514
rect 11683 20968 12053 21341
rect 11526 20958 11683 20968
rect 12043 15122 12053 20968
rect 12227 20805 12237 21700
rect 12820 21739 14370 21859
rect 12468 21521 12478 21585
rect 12678 21521 12688 21585
rect 12820 21063 12940 21739
rect 13511 21508 13521 21556
rect 13285 21408 13295 21508
rect 13347 21456 13521 21508
rect 13573 21456 13583 21556
rect 13656 21456 13666 21556
rect 13718 21508 13728 21556
rect 13718 21456 13866 21508
rect 13347 21408 13357 21456
rect 13856 21408 13866 21456
rect 13918 21408 13928 21508
rect 14250 21447 14370 21739
rect 14984 21579 14994 21656
rect 14525 21527 14535 21579
rect 14735 21527 14994 21579
rect 14248 21395 14258 21447
rect 14358 21395 14370 21447
rect 13044 21267 13054 21323
rect 13254 21267 13264 21323
rect 14250 21321 14370 21395
rect 13511 21198 13521 21298
rect 13573 21250 13583 21298
rect 14250 21269 14260 21321
rect 14360 21269 14370 21321
rect 13573 21198 13866 21250
rect 13856 21066 13866 21198
rect 13918 21066 13928 21250
rect 12820 21011 12830 21063
rect 12930 21011 12940 21063
rect 12820 20934 12940 21011
rect 13656 20992 13666 21040
rect 12819 20882 12824 20934
rect 12929 20882 12940 20934
rect 13285 20892 13295 20992
rect 13347 20940 13666 20992
rect 13718 20940 13728 21040
rect 13347 20892 13357 20940
rect 12227 20753 12478 20805
rect 12678 20753 12688 20805
rect 12227 19256 12237 20753
rect 12820 20672 12940 20882
rect 13949 20747 13959 20811
rect 14159 20747 14169 20811
rect 12817 20620 12827 20672
rect 12927 20620 12940 20672
rect 12820 20547 12940 20620
rect 12820 20495 12830 20547
rect 12930 20495 12940 20547
rect 12468 19973 12478 20037
rect 12678 19973 12688 20037
rect 12820 19515 12940 20495
rect 13511 20476 13521 20524
rect 13285 20351 13295 20476
rect 13347 20424 13521 20476
rect 13573 20424 13583 20524
rect 13347 20351 13357 20424
rect 13044 20235 13054 20291
rect 13254 20235 13264 20291
rect 14250 20289 14370 21269
rect 14525 21009 14535 21065
rect 14735 21009 14745 21065
rect 14525 20493 14535 20549
rect 14735 20493 14745 20549
rect 13656 20166 13666 20266
rect 13718 20218 13728 20266
rect 14250 20237 14260 20289
rect 14360 20237 14370 20289
rect 13718 20166 13866 20218
rect 13856 20118 13866 20166
rect 13918 20118 13928 20218
rect 14250 20155 14370 20237
rect 14250 20103 14260 20155
rect 14360 20103 14370 20155
rect 14250 19900 14370 20103
rect 14984 20031 14994 21527
rect 14525 19979 14535 20031
rect 14735 19979 14994 20031
rect 14250 19848 14262 19900
rect 14362 19848 14372 19900
rect 13044 19719 13054 19775
rect 13254 19719 13264 19775
rect 14250 19773 14370 19848
rect 13511 19650 13521 19750
rect 13573 19702 13583 19750
rect 14250 19721 14260 19773
rect 14360 19721 14370 19773
rect 13573 19650 13866 19702
rect 13856 19518 13866 19650
rect 13918 19518 13928 19702
rect 12820 19463 12830 19515
rect 12930 19463 12940 19515
rect 12820 19381 12940 19463
rect 13656 19444 13666 19492
rect 12819 19329 12829 19381
rect 12929 19329 12940 19381
rect 13285 19344 13295 19444
rect 13347 19392 13666 19444
rect 13718 19392 13728 19492
rect 13347 19344 13357 19392
rect 12227 19204 12478 19256
rect 12678 19204 12688 19256
rect 12227 17709 12237 19204
rect 12820 19129 12940 19329
rect 13949 19199 13959 19263
rect 14159 19199 14169 19263
rect 12820 19077 12832 19129
rect 12932 19077 12942 19129
rect 12820 18999 12940 19077
rect 12820 18947 12830 18999
rect 12930 18947 12940 18999
rect 12468 18425 12478 18489
rect 12678 18425 12688 18489
rect 12820 17967 12940 18947
rect 13511 18928 13521 18976
rect 13285 18802 13295 18928
rect 13347 18876 13521 18928
rect 13573 18876 13583 18976
rect 13347 18802 13357 18876
rect 13044 18687 13054 18743
rect 13254 18687 13264 18743
rect 14250 18741 14370 19721
rect 14525 19461 14535 19517
rect 14735 19461 14745 19517
rect 14525 18945 14535 19001
rect 14735 18945 14745 19001
rect 13656 18618 13666 18718
rect 13718 18670 13728 18718
rect 14249 18689 14259 18741
rect 14359 18689 14370 18741
rect 13718 18618 13866 18670
rect 13856 18570 13866 18618
rect 13918 18570 13928 18670
rect 14250 18604 14370 18689
rect 14250 18552 14262 18604
rect 14362 18552 14372 18604
rect 14250 18342 14370 18552
rect 14984 18483 14994 19979
rect 14525 18431 14535 18483
rect 14735 18431 14994 18483
rect 14250 18290 14260 18342
rect 14360 18290 14370 18342
rect 13044 18171 13054 18227
rect 13254 18171 13264 18227
rect 14250 18225 14370 18290
rect 13511 18102 13521 18202
rect 13573 18154 13583 18202
rect 14250 18173 14260 18225
rect 14360 18173 14370 18225
rect 13573 18102 13866 18154
rect 13856 17970 13866 18102
rect 13918 17970 13928 18154
rect 12820 17915 12830 17967
rect 12930 17915 12940 17967
rect 12820 17836 12940 17915
rect 13656 17896 13666 17944
rect 12820 17784 12831 17836
rect 12931 17784 12941 17836
rect 13285 17796 13295 17896
rect 13347 17844 13666 17896
rect 13718 17844 13728 17944
rect 13347 17796 13357 17844
rect 12227 17657 12478 17709
rect 12678 17657 12688 17709
rect 12227 16161 12237 17657
rect 12820 17574 12940 17784
rect 13949 17651 13959 17715
rect 14159 17651 14169 17715
rect 12819 17522 12829 17574
rect 12929 17522 12940 17574
rect 12820 17451 12940 17522
rect 12820 17399 12830 17451
rect 12930 17399 12940 17451
rect 12468 16877 12478 16941
rect 12678 16877 12688 16941
rect 12820 16419 12940 17399
rect 13511 17380 13521 17428
rect 13285 17254 13295 17380
rect 13347 17328 13521 17380
rect 13573 17328 13583 17428
rect 13347 17254 13357 17328
rect 13285 17248 13357 17254
rect 13044 17139 13054 17195
rect 13254 17139 13264 17195
rect 14250 17193 14370 18173
rect 14525 17913 14535 17969
rect 14735 17913 14745 17969
rect 14525 17397 14535 17453
rect 14735 17397 14745 17453
rect 13656 17070 13666 17170
rect 13718 17122 13728 17170
rect 14250 17141 14260 17193
rect 14360 17141 14370 17193
rect 13718 17070 13866 17122
rect 13856 17022 13866 17070
rect 13918 17022 13928 17122
rect 14250 17056 14370 17141
rect 14248 17004 14258 17056
rect 14358 17004 14370 17056
rect 14250 16800 14370 17004
rect 14984 16935 14994 18431
rect 14525 16883 14535 16935
rect 14735 16883 14994 16935
rect 14249 16748 14259 16800
rect 14359 16748 14370 16800
rect 13044 16623 13054 16679
rect 13254 16623 13264 16679
rect 14250 16677 14370 16748
rect 13511 16554 13521 16654
rect 13573 16606 13583 16654
rect 14250 16625 14260 16677
rect 14360 16625 14370 16677
rect 13573 16554 13866 16606
rect 12820 16367 12830 16419
rect 12930 16367 12940 16419
rect 13856 16406 13866 16554
rect 13918 16406 13928 16606
rect 12820 16292 12940 16367
rect 13656 16348 13666 16396
rect 12820 16240 12830 16292
rect 12930 16240 12940 16292
rect 13285 16248 13295 16348
rect 13347 16296 13666 16348
rect 13718 16296 13728 16396
rect 13347 16248 13357 16296
rect 12227 16109 12478 16161
rect 12678 16109 12688 16161
rect 12227 15179 12237 16109
rect 12820 16027 12940 16240
rect 13949 16103 13959 16167
rect 14159 16103 14169 16167
rect 12820 15975 12830 16027
rect 12930 15975 12940 16027
rect 12820 15903 12940 15975
rect 12820 15851 12830 15903
rect 12930 15851 12940 15903
rect 13511 15832 13521 15880
rect 13285 15732 13295 15832
rect 13347 15780 13521 15832
rect 13573 15780 13583 15880
rect 13347 15732 13357 15780
rect 13044 15591 13054 15647
rect 13254 15591 13264 15647
rect 14250 15645 14370 16625
rect 14525 16365 14535 16421
rect 14735 16365 14745 16421
rect 14524 15849 14534 15905
rect 14734 15849 14744 15905
rect 13656 15522 13666 15622
rect 13718 15574 13728 15622
rect 14250 15593 14260 15645
rect 14360 15593 14370 15645
rect 13718 15522 13866 15574
rect 13856 15474 13866 15522
rect 13918 15474 13928 15574
rect 14250 15522 14370 15593
rect 14250 15470 14262 15522
rect 14362 15470 14372 15522
rect 14250 15446 14370 15470
rect 12468 15329 12478 15393
rect 12678 15329 12688 15393
rect 14984 15387 14994 16883
rect 14525 15335 14535 15387
rect 14735 15335 14994 15387
rect 14984 15315 14994 15335
rect 15106 16340 15116 21656
rect 15726 17060 15736 22467
rect 15927 17060 15937 22467
rect 16576 22449 16676 22578
rect 16576 22397 16883 22449
rect 17006 22397 17016 22449
rect 16576 22384 16676 22397
rect 16086 22332 16096 22384
rect 16156 22332 16212 22384
rect 16272 22332 16676 22384
rect 16086 21868 16166 22332
rect 16086 21816 16096 21868
rect 16156 21816 16166 21868
rect 16086 21352 16166 21816
rect 16202 22074 16212 22126
rect 16272 22074 16282 22126
rect 16202 21868 16282 22074
rect 17314 21991 17324 22497
rect 16926 21939 16936 21991
rect 17059 21939 17324 21991
rect 16202 21816 16883 21868
rect 17006 21816 17015 21868
rect 16202 21610 16282 21816
rect 16202 21558 16212 21610
rect 16272 21558 16282 21610
rect 17314 21410 17324 21939
rect 16925 21358 16935 21410
rect 17059 21358 17324 21410
rect 16086 21300 16096 21352
rect 16156 21300 16166 21352
rect 17314 21143 17324 21358
rect 17475 21143 17485 22497
rect 16086 21042 16096 21094
rect 16156 21042 16166 21094
rect 16086 20578 16166 21042
rect 16086 20526 16096 20578
rect 16156 20526 16166 20578
rect 16086 20062 16166 20526
rect 16202 20784 16212 20836
rect 16272 20784 16282 20836
rect 16202 20578 16282 20784
rect 16202 20526 16883 20578
rect 16996 20526 17006 20578
rect 16202 20320 16282 20526
rect 16202 20268 16212 20320
rect 16272 20268 16282 20320
rect 17320 20120 17330 21143
rect 16926 20068 16936 20120
rect 17059 20068 17330 20120
rect 16086 20010 16096 20062
rect 16156 20010 16166 20062
rect 16086 19752 16096 19804
rect 16156 19752 16166 19804
rect 16086 19288 16166 19752
rect 16086 19236 16096 19288
rect 16156 19236 16166 19288
rect 16086 18778 16166 19236
rect 16202 19494 16212 19546
rect 16272 19494 16282 19546
rect 16202 19288 16282 19494
rect 16202 19236 16883 19288
rect 16996 19236 17006 19288
rect 16202 19030 16282 19236
rect 16202 18978 16212 19030
rect 16272 18978 16282 19030
rect 17320 18830 17330 20068
rect 16926 18778 16936 18830
rect 17059 18778 17330 18830
rect 16086 18714 16096 18778
rect 16160 18714 16170 18778
rect 16086 18462 16096 18514
rect 16156 18462 16166 18514
rect 16086 17998 16166 18462
rect 16086 17946 16096 17998
rect 16156 17946 16166 17998
rect 16086 17482 16166 17946
rect 16202 18204 16212 18256
rect 16272 18204 16282 18256
rect 16202 17998 16282 18204
rect 16202 17946 16883 17998
rect 16996 17946 17006 17998
rect 16202 17740 16282 17946
rect 16202 17688 16212 17740
rect 16272 17688 16282 17740
rect 17320 17540 17330 18778
rect 16926 17488 16936 17540
rect 17059 17490 17330 17540
rect 17469 18131 17479 21143
rect 20371 18779 20450 25496
rect 20762 25493 20797 25500
rect 20762 25490 25207 25493
rect 20797 25483 25207 25490
rect 22120 25360 24248 25370
rect 22178 25247 24248 25257
rect 22694 25092 22746 25093
rect 23610 25092 23662 25093
rect 22694 25083 24542 25092
rect 22746 24992 23610 25083
rect 22694 24913 22746 24923
rect 23662 24992 24542 25083
rect 23132 24912 23226 24922
rect 23610 24913 23662 24923
rect 23132 24765 23226 24775
rect 22120 24709 22178 24719
rect 22213 24654 22307 24664
rect 22213 24507 22307 24517
rect 24048 24654 24142 24664
rect 24048 24507 24142 24517
rect 22475 24466 22675 24476
rect 22475 24404 22675 24414
rect 22933 24466 23133 24476
rect 22933 24404 23133 24414
rect 23391 24466 23591 24476
rect 23391 24404 23591 24414
rect 23849 24466 24049 24476
rect 23849 24404 24049 24414
rect 20736 24342 20819 24352
rect 20736 24232 20819 24242
rect 22575 24342 22675 24404
rect 22575 24232 22675 24242
rect 22765 24342 22865 24352
rect 20726 24156 20839 24166
rect 20726 24046 20839 24056
rect 22307 24156 22407 24166
rect 22307 23979 22407 24056
rect 22765 23979 22865 24242
rect 23033 24156 23133 24404
rect 23033 24046 23133 24056
rect 23223 24342 23323 24352
rect 23223 23979 23323 24242
rect 23491 24156 23591 24404
rect 23949 24342 24049 24404
rect 23949 24232 24049 24242
rect 23491 24046 23591 24056
rect 23681 24156 23781 24166
rect 23681 23979 23781 24056
rect 22307 23969 22507 23979
rect 22307 23907 22507 23917
rect 22765 23969 22965 23979
rect 22765 23907 22965 23917
rect 23223 23969 23423 23979
rect 23223 23907 23423 23917
rect 23681 23969 23881 23979
rect 23681 23907 23881 23917
rect 22214 23865 22308 23875
rect 22214 23718 22308 23728
rect 24046 23865 24140 23875
rect 24046 23718 24140 23728
rect 22111 23683 22185 23693
rect 21347 23600 21659 23610
rect 21659 23382 22111 23600
rect 21347 23372 21659 23382
rect 22066 23052 22111 23062
rect 23131 23654 23225 23664
rect 23131 23507 23225 23517
rect 22694 23460 22746 23470
rect 23610 23460 23662 23470
rect 22746 23300 23610 23393
rect 24442 23393 24542 24992
rect 25311 24965 25792 24975
rect 25311 24833 25384 24965
rect 25436 24833 25740 24965
rect 25384 24755 25436 24765
rect 25740 24755 25792 24765
rect 25207 24324 25311 24334
rect 25512 24669 25564 24679
rect 25512 24083 25564 24469
rect 25512 23994 25564 24004
rect 25868 24669 25920 24679
rect 25868 24249 25920 24469
rect 29707 24249 29886 24259
rect 25868 24069 29707 24249
rect 25868 23960 25920 24069
rect 25868 23879 25920 23889
rect 25424 23855 25476 23865
rect 25424 23510 25476 23784
rect 25780 23855 25832 23865
rect 25780 23510 25832 23784
rect 23662 23300 24542 23393
rect 22694 23293 24542 23300
rect 24611 23500 25989 23510
rect 22694 23290 22746 23293
rect 23610 23290 23741 23293
rect 22185 23055 22293 23062
rect 22185 23052 23409 23055
rect 22293 23045 23409 23052
rect 22024 21625 22066 21899
rect 22404 22865 23409 22875
rect 23619 22776 23741 23290
rect 24611 23218 25989 23228
rect 24701 23018 24842 23028
rect 24842 23008 25109 23018
rect 26151 23017 26223 24069
rect 29707 24058 29886 24068
rect 24842 22956 24907 23008
rect 24701 22946 24842 22956
rect 24907 22946 25109 22956
rect 25741 23007 26223 23017
rect 25943 22955 26223 23007
rect 25741 22945 26223 22955
rect 23955 22917 24166 22927
rect 23333 22766 23742 22776
rect 23333 22691 23742 22701
rect 22571 22673 22627 22683
rect 22571 22523 22627 22533
rect 22404 22407 23166 22417
rect 22404 22343 22666 22407
rect 22404 22333 23166 22343
rect 23619 22060 23741 22691
rect 23333 22050 23742 22060
rect 23333 21975 23742 21985
rect 22404 21866 23955 21876
rect 22293 21625 23955 21627
rect 22024 21617 23955 21625
rect 22024 21615 22293 21617
rect 22024 21614 22184 21615
rect 23955 21606 24166 21616
rect 20371 18703 20450 18713
rect 30362 20775 30542 20785
rect 18099 18131 18521 18141
rect 17469 17743 18099 18131
rect 17469 17490 17479 17743
rect 18099 17733 18521 17743
rect 30362 17647 30542 20632
rect 17059 17488 17479 17490
rect 16086 17430 16096 17482
rect 16156 17430 16166 17482
rect 15726 16967 15937 17060
rect 16086 17172 16096 17224
rect 16156 17172 16166 17224
rect 16086 16806 16166 17172
rect 17320 17029 17479 17488
rect 30358 17477 30367 17647
rect 30537 17477 30546 17647
rect 30362 17472 30542 17477
rect 17320 17028 17429 17029
rect 16873 16852 16883 16916
rect 17023 16852 17033 16916
rect 15364 16726 15374 16806
rect 15447 16726 16166 16806
rect 17206 16652 17216 17028
rect 16909 16600 16919 16652
rect 17059 16600 17216 16652
rect 15106 16316 16507 16340
rect 16873 16336 16883 16400
rect 17023 16336 17033 16400
rect 15106 16208 15334 16316
rect 16377 16208 16507 16316
rect 15106 16186 16507 16208
rect 15106 15834 15116 16186
rect 16317 16083 16507 16186
rect 15570 15941 15580 16015
rect 16180 15941 16190 16015
rect 15106 15315 15155 15834
rect 14984 15307 15155 15315
rect 15251 15307 15261 15834
rect 16317 15307 16344 16083
rect 14984 15302 15261 15307
rect 14984 15179 15038 15302
rect 12227 15125 12309 15179
rect 12461 15125 13299 15179
rect 13447 15125 15038 15179
rect 15755 15281 16344 15307
rect 15755 15161 15767 15281
rect 16246 15258 16344 15281
rect 16492 15258 16507 16083
rect 16753 15749 16763 16108
rect 16828 15749 16838 16108
rect 17206 16042 17216 16600
rect 17351 16042 17429 17028
rect 17208 15727 17218 16042
rect 16873 15675 16883 15727
rect 16959 15675 17218 15727
rect 16753 15295 16763 15654
rect 16828 15295 16838 15654
rect 17208 15467 17218 15675
rect 17189 15415 17218 15467
rect 16246 15161 16507 15258
rect 15755 15146 16507 15161
rect 12227 15122 12237 15125
rect 12043 15010 12237 15122
rect 17208 15049 17218 15415
rect 17350 15050 17429 16042
rect 17577 15050 17587 17029
rect 17350 15049 17587 15050
rect 17274 15048 17587 15049
rect 17423 14978 17587 15048
rect 30362 13028 30542 13038
rect 13963 12273 14168 12283
rect 7845 11892 13963 12273
rect 1903 10420 2303 10430
rect 2678 10420 2872 10559
rect 7845 10480 8226 11892
rect 13963 11882 14168 11892
rect 25902 11405 26136 11414
rect 17726 11404 26136 11405
rect 17726 11104 25902 11404
rect 17726 11015 17910 11104
rect 25708 11015 25902 11104
rect 17726 11005 25902 11015
rect 2303 10407 2872 10420
rect 2303 10020 2688 10407
rect 1903 10010 2303 10020
rect 2678 3829 2688 10020
rect 2862 10404 2872 10407
rect 2862 10350 2944 10404
rect 3096 10350 3934 10404
rect 4082 10350 5673 10404
rect 2862 9420 2872 10350
rect 5619 10227 5673 10350
rect 6390 10368 7142 10383
rect 6390 10248 6402 10368
rect 6881 10271 7142 10368
rect 6881 10248 6979 10271
rect 5619 10222 5896 10227
rect 6390 10222 6979 10248
rect 5619 10214 5790 10222
rect 3103 10136 3113 10200
rect 3313 10136 3323 10200
rect 5619 10194 5629 10214
rect 5160 10142 5170 10194
rect 5370 10142 5629 10194
rect 4885 10059 5005 10083
rect 4491 10007 4501 10055
rect 3679 9882 3689 9938
rect 3889 9882 3899 9938
rect 4291 9907 4301 10007
rect 4353 9955 4501 10007
rect 4553 9955 4563 10055
rect 4885 10007 4897 10059
rect 4997 10007 5007 10059
rect 4353 9907 4363 9955
rect 4885 9936 5005 10007
rect 4885 9884 4895 9936
rect 4995 9884 5005 9936
rect 3920 9697 3930 9797
rect 3982 9749 3992 9797
rect 3982 9697 4156 9749
rect 3455 9626 3465 9678
rect 3565 9626 3575 9678
rect 4146 9649 4156 9697
rect 4208 9649 4218 9749
rect 3455 9554 3575 9626
rect 3455 9502 3465 9554
rect 3565 9502 3575 9554
rect 2862 9368 3113 9420
rect 3313 9368 3323 9420
rect 2862 7872 2872 9368
rect 3455 9289 3575 9502
rect 4584 9362 4594 9426
rect 4794 9362 4804 9426
rect 3455 9237 3465 9289
rect 3565 9237 3575 9289
rect 3455 9162 3575 9237
rect 3920 9181 3930 9281
rect 3982 9233 3992 9281
rect 3982 9181 4301 9233
rect 3455 9110 3465 9162
rect 3565 9110 3575 9162
rect 4291 9133 4301 9181
rect 4353 9133 4363 9233
rect 3103 8588 3113 8652
rect 3313 8588 3323 8652
rect 3455 8130 3575 9110
rect 4491 8975 4501 9123
rect 3679 8850 3689 8906
rect 3889 8850 3899 8906
rect 4146 8875 4156 8975
rect 4208 8923 4501 8975
rect 4553 8923 4563 9123
rect 4208 8875 4218 8923
rect 4885 8904 5005 9884
rect 5159 9624 5169 9680
rect 5369 9624 5379 9680
rect 5160 9108 5170 9164
rect 5370 9108 5380 9164
rect 4885 8852 4895 8904
rect 4995 8852 5005 8904
rect 4885 8781 5005 8852
rect 4884 8729 4894 8781
rect 4994 8729 5005 8781
rect 4885 8525 5005 8729
rect 5619 8646 5629 10142
rect 5160 8594 5170 8646
rect 5370 8594 5629 8646
rect 4491 8459 4501 8507
rect 3679 8334 3689 8390
rect 3889 8334 3899 8390
rect 4291 8359 4301 8459
rect 4353 8407 4501 8459
rect 4553 8407 4563 8507
rect 4883 8473 4893 8525
rect 4993 8473 5005 8525
rect 4353 8359 4363 8407
rect 4885 8388 5005 8473
rect 4885 8336 4895 8388
rect 4995 8336 5005 8388
rect 3920 8275 3992 8281
rect 3920 8149 3930 8275
rect 3982 8201 3992 8275
rect 3982 8149 4156 8201
rect 3455 8078 3465 8130
rect 3565 8078 3575 8130
rect 4146 8101 4156 8149
rect 4208 8101 4218 8201
rect 3455 8007 3575 8078
rect 3454 7955 3464 8007
rect 3564 7955 3575 8007
rect 2862 7820 3113 7872
rect 3313 7820 3323 7872
rect 2862 6325 2872 7820
rect 3455 7745 3575 7955
rect 4584 7814 4594 7878
rect 4794 7814 4804 7878
rect 3455 7693 3466 7745
rect 3566 7693 3576 7745
rect 3455 7614 3575 7693
rect 3920 7633 3930 7733
rect 3982 7685 3992 7733
rect 3982 7633 4301 7685
rect 3455 7562 3465 7614
rect 3565 7562 3575 7614
rect 4291 7585 4301 7633
rect 4353 7585 4363 7685
rect 3103 7040 3113 7104
rect 3313 7040 3323 7104
rect 3455 6582 3575 7562
rect 4491 7427 4501 7559
rect 3679 7302 3689 7358
rect 3889 7302 3899 7358
rect 4146 7327 4156 7427
rect 4208 7375 4501 7427
rect 4553 7375 4563 7559
rect 4208 7327 4218 7375
rect 4885 7356 5005 8336
rect 5160 8076 5170 8132
rect 5370 8076 5380 8132
rect 5160 7560 5170 7616
rect 5370 7560 5380 7616
rect 4885 7304 4895 7356
rect 4995 7304 5005 7356
rect 4885 7239 5005 7304
rect 4885 7187 4895 7239
rect 4995 7187 5005 7239
rect 4885 6977 5005 7187
rect 5619 7098 5629 8594
rect 5160 7046 5170 7098
rect 5370 7046 5629 7098
rect 4491 6911 4501 6959
rect 3679 6786 3689 6842
rect 3889 6786 3899 6842
rect 4291 6811 4301 6911
rect 4353 6859 4501 6911
rect 4553 6859 4563 6959
rect 4885 6925 4897 6977
rect 4997 6925 5007 6977
rect 4353 6811 4363 6859
rect 4885 6840 5005 6925
rect 4884 6788 4894 6840
rect 4994 6788 5005 6840
rect 3920 6601 3930 6727
rect 3982 6653 3992 6727
rect 3982 6601 4156 6653
rect 3455 6530 3465 6582
rect 3565 6530 3575 6582
rect 4146 6553 4156 6601
rect 4208 6553 4218 6653
rect 3455 6452 3575 6530
rect 3455 6400 3467 6452
rect 3567 6400 3577 6452
rect 2862 6273 3113 6325
rect 3313 6273 3323 6325
rect 2862 4776 2872 6273
rect 3455 6200 3575 6400
rect 4584 6266 4594 6330
rect 4794 6266 4804 6330
rect 3454 6148 3464 6200
rect 3564 6148 3575 6200
rect 3455 6066 3575 6148
rect 3920 6085 3930 6185
rect 3982 6137 3992 6185
rect 3982 6085 4301 6137
rect 3455 6014 3465 6066
rect 3565 6014 3575 6066
rect 4291 6037 4301 6085
rect 4353 6037 4363 6137
rect 3103 5492 3113 5556
rect 3313 5492 3323 5556
rect 3455 5034 3575 6014
rect 4491 5879 4501 6011
rect 3679 5754 3689 5810
rect 3889 5754 3899 5810
rect 4146 5779 4156 5879
rect 4208 5827 4501 5879
rect 4553 5827 4563 6011
rect 4208 5779 4218 5827
rect 4885 5808 5005 6788
rect 5160 6528 5170 6584
rect 5370 6528 5380 6584
rect 5160 6012 5170 6068
rect 5370 6012 5380 6068
rect 4885 5756 4895 5808
rect 4995 5756 5005 5808
rect 4885 5681 5005 5756
rect 4885 5629 4897 5681
rect 4997 5629 5007 5681
rect 4885 5426 5005 5629
rect 5619 5550 5629 7046
rect 5160 5498 5170 5550
rect 5370 5498 5629 5550
rect 4491 5363 4501 5411
rect 3679 5238 3689 5294
rect 3889 5238 3899 5294
rect 4291 5263 4301 5363
rect 4353 5311 4501 5363
rect 4553 5311 4563 5411
rect 4885 5374 4895 5426
rect 4995 5374 5005 5426
rect 4353 5263 4363 5311
rect 4885 5292 5005 5374
rect 4885 5240 4895 5292
rect 4995 5240 5005 5292
rect 3920 5053 3930 5178
rect 3982 5105 3992 5178
rect 3982 5053 4156 5105
rect 3455 4982 3465 5034
rect 3565 4982 3575 5034
rect 4146 5005 4156 5053
rect 4208 5005 4218 5105
rect 3455 4909 3575 4982
rect 3452 4857 3462 4909
rect 3562 4857 3575 4909
rect 2862 4724 3113 4776
rect 3313 4724 3323 4776
rect 2862 3829 2872 4724
rect 3455 4647 3575 4857
rect 4584 4718 4594 4782
rect 4794 4718 4804 4782
rect 3454 4595 3459 4647
rect 3564 4595 3575 4647
rect 3455 4518 3575 4595
rect 3920 4537 3930 4637
rect 3982 4589 3992 4637
rect 3982 4537 4301 4589
rect 3455 4466 3465 4518
rect 3565 4466 3575 4518
rect 4291 4489 4301 4537
rect 4353 4489 4363 4589
rect 3103 3944 3113 4008
rect 3313 3944 3323 4008
rect 3455 3790 3575 4466
rect 4491 4331 4501 4463
rect 3679 4206 3689 4262
rect 3889 4206 3899 4262
rect 4146 4231 4156 4331
rect 4208 4279 4501 4331
rect 4553 4279 4563 4463
rect 4208 4231 4218 4279
rect 4885 4260 5005 5240
rect 5160 4980 5170 5036
rect 5370 4980 5380 5036
rect 5160 4464 5170 4520
rect 5370 4464 5380 4520
rect 4885 4208 4895 4260
rect 4995 4208 5005 4260
rect 4885 4134 5005 4208
rect 3920 4021 3930 4121
rect 3982 4073 3992 4121
rect 4491 4073 4501 4121
rect 3982 4021 4156 4073
rect 4146 3973 4156 4021
rect 4208 3973 4218 4073
rect 4291 3973 4301 4073
rect 4353 4021 4501 4073
rect 4553 4021 4563 4121
rect 4883 4082 4893 4134
rect 4993 4082 5005 4134
rect 4353 3973 4363 4021
rect 4885 3790 5005 4082
rect 5619 4002 5629 5498
rect 5160 3950 5170 4002
rect 5370 3950 5629 4002
rect 5619 3873 5629 3950
rect 5741 9695 5790 10214
rect 5886 9695 5896 10222
rect 5741 9343 5751 9695
rect 6205 9514 6215 9588
rect 6815 9514 6825 9588
rect 6952 9446 6979 10222
rect 7127 9446 7142 10271
rect 7388 9875 7398 10234
rect 7463 9875 7473 10234
rect 7843 10114 7853 10480
rect 7824 10062 7853 10114
rect 7843 9854 7853 10062
rect 7508 9802 7518 9854
rect 7594 9802 7853 9854
rect 6952 9343 7142 9446
rect 7388 9421 7398 9780
rect 7463 9421 7473 9780
rect 7843 9487 7853 9802
rect 7985 10479 8226 10480
rect 7985 9487 8064 10479
rect 5741 9321 7142 9343
rect 5741 9213 5969 9321
rect 7012 9213 7142 9321
rect 5741 9189 7142 9213
rect 5741 3873 5751 9189
rect 7508 9129 7518 9193
rect 7658 9129 7668 9193
rect 7841 8929 7851 9487
rect 7544 8877 7554 8929
rect 7694 8877 7851 8929
rect 5987 8666 5997 8746
rect 6082 8666 6801 8746
rect 6361 8370 6572 8463
rect 3455 3670 5005 3790
rect 6361 2963 6371 8370
rect 6562 2963 6572 8370
rect 6721 8258 6801 8666
rect 7508 8613 7518 8677
rect 7658 8613 7668 8677
rect 7841 8501 7851 8877
rect 7986 8501 8064 9487
rect 6721 8206 6731 8258
rect 6791 8206 6801 8258
rect 7954 8500 8064 8501
rect 8212 10380 8226 10479
rect 21823 10654 21877 11005
rect 25902 10994 26136 11004
rect 8212 8500 8222 10380
rect 18132 10135 18218 10178
rect 18132 9830 18142 10135
rect 18132 9462 18218 9830
rect 21823 10166 21877 10318
rect 21823 9820 21877 9830
rect 25483 10125 25569 10178
rect 25559 9830 25569 10125
rect 18132 9452 18451 9462
rect 18132 9368 18142 9452
rect 18132 9358 18451 9368
rect 18950 9444 19311 9459
rect 19299 9377 19311 9444
rect 18950 9359 19311 9377
rect 24014 9441 24379 9459
rect 24363 9374 24379 9441
rect 24014 9359 24379 9374
rect 7954 8042 8115 8500
rect 6721 7948 6731 8000
rect 6791 7948 6801 8000
rect 6721 7484 6801 7948
rect 7955 7942 8114 8042
rect 7561 7890 7571 7942
rect 7694 7940 8114 7942
rect 7694 7890 7965 7940
rect 6721 7432 6731 7484
rect 6791 7432 6801 7484
rect 6721 6968 6801 7432
rect 6837 7690 6847 7742
rect 6907 7690 6917 7742
rect 6837 7484 6917 7690
rect 6837 7432 7518 7484
rect 7631 7432 7641 7484
rect 6837 7226 6917 7432
rect 6837 7174 6847 7226
rect 6907 7174 6917 7226
rect 6721 6916 6731 6968
rect 6791 6916 6801 6968
rect 6721 6658 6731 6710
rect 6791 6658 6801 6710
rect 6721 6194 6801 6658
rect 7955 6652 7965 7890
rect 7561 6600 7571 6652
rect 7694 6600 7965 6652
rect 6721 6142 6731 6194
rect 6791 6142 6801 6194
rect 6721 5678 6801 6142
rect 6837 6400 6847 6452
rect 6907 6400 6917 6452
rect 6837 6194 6917 6400
rect 6837 6142 7518 6194
rect 7631 6142 7641 6194
rect 6837 5936 6917 6142
rect 6837 5884 6847 5936
rect 6907 5884 6917 5936
rect 6721 5626 6731 5678
rect 6791 5626 6801 5678
rect 6721 5368 6731 5420
rect 6791 5368 6801 5420
rect 6721 4904 6801 5368
rect 7955 5362 7965 6600
rect 7561 5310 7571 5362
rect 7694 5310 7965 5362
rect 6721 4852 6731 4904
rect 6791 4852 6801 4904
rect 6721 4388 6801 4852
rect 6837 5110 6847 5162
rect 6907 5110 6917 5162
rect 6837 4904 6917 5110
rect 6837 4852 7518 4904
rect 7631 4852 7641 4904
rect 6837 4646 6917 4852
rect 6837 4594 6847 4646
rect 6907 4594 6917 4646
rect 6721 4336 6731 4388
rect 6791 4336 6801 4388
rect 7955 4287 7965 5310
rect 8104 4287 8114 7940
rect 18058 7296 18634 7306
rect 18058 7221 18634 7231
rect 18676 7047 18728 7048
rect 18673 7038 18731 7047
rect 18673 7037 18676 7038
rect 18728 7037 18731 7038
rect 11501 6554 11886 6563
rect 18673 6229 18731 6239
rect 19225 6917 19311 9359
rect 19341 9254 19727 9274
rect 19341 9187 19377 9254
rect 19726 9187 19727 9254
rect 19341 9174 19727 9187
rect 19341 8782 19427 9174
rect 19341 8204 19427 8214
rect 24293 8782 24379 9359
rect 25483 9274 25569 9830
rect 26498 9459 26678 9469
rect 26498 9288 26678 9298
rect 24293 8204 24379 8214
rect 24409 9258 24783 9274
rect 24409 9191 24434 9258
rect 24409 9174 24783 9191
rect 25148 9258 25569 9274
rect 25538 9188 25569 9258
rect 25148 9174 25569 9188
rect 21831 7970 21887 7980
rect 21831 7618 21887 7628
rect 19451 7568 19661 7578
rect 19451 7450 19661 7511
rect 24063 7568 24273 7578
rect 19451 7393 19474 7450
rect 19451 7383 19661 7393
rect 21904 7454 22114 7466
rect 22105 7390 22114 7454
rect 21604 7135 21814 7145
rect 21604 7003 21814 7078
rect 21604 6936 21814 6946
rect 21904 7002 22114 7390
rect 24063 7137 24273 7511
rect 24063 7070 24273 7080
rect 21904 6935 22114 6945
rect 24409 6917 24495 9174
rect 30362 8230 30542 12891
rect 30362 8077 30542 8087
rect 19225 6907 19426 6917
rect 11501 5732 11886 6169
rect 19225 5835 19274 6907
rect 24291 6907 24495 6917
rect 21830 6886 21888 6896
rect 21830 6537 21888 6547
rect 19426 5835 19428 6343
rect 19225 5766 19428 5835
rect 24443 5835 24495 6907
rect 24291 5825 24495 5835
rect 17724 5732 18506 5733
rect 11501 5667 18506 5732
rect 11501 5573 17832 5667
rect 18385 5573 18506 5667
rect 19446 5691 19926 5701
rect 19446 5623 19926 5633
rect 21904 5693 22384 5703
rect 21904 5625 22384 5635
rect 11501 5442 18506 5573
rect 11501 5432 24768 5442
rect 11501 5347 17834 5432
rect 17447 5343 17834 5347
rect 17447 5333 24768 5343
rect 17447 5332 17727 5333
rect 6721 4078 6731 4130
rect 6791 4078 6801 4130
rect 6721 3614 6801 4078
rect 7949 4072 7959 4287
rect 7560 4020 7570 4072
rect 7694 4020 7959 4072
rect 6721 3562 6731 3614
rect 6791 3562 6801 3614
rect 6721 3098 6801 3562
rect 6837 3820 6847 3872
rect 6907 3820 6917 3872
rect 6837 3614 6917 3820
rect 6837 3562 7518 3614
rect 7641 3562 7650 3614
rect 6837 3356 6917 3562
rect 7949 3491 7959 4020
rect 7561 3439 7571 3491
rect 7694 3439 7959 3491
rect 6837 3304 6847 3356
rect 6907 3304 6917 3356
rect 6721 3046 6731 3098
rect 6791 3046 6847 3098
rect 6907 3046 7358 3098
rect 7178 3033 7358 3046
rect 7178 2981 7518 3033
rect 7641 2981 7651 3033
rect 7178 2767 7358 2981
rect 7949 2933 7959 3439
rect 8110 2933 8120 4287
rect 7178 2648 7358 2658
<< via2 >>
rect 11865 32876 14344 32983
rect 10935 30961 11665 31121
rect 3549 27072 4125 27082
rect 3549 27017 4125 27072
rect 4164 26025 4167 26823
rect 4167 26025 4219 26823
rect 4219 26025 4222 26823
rect 12999 30777 13063 31777
rect 12122 29540 12186 30540
rect 13875 29540 13939 30540
rect 7322 27743 7378 27756
rect 7322 27424 7326 27743
rect 7326 27424 7378 27743
rect 7322 27414 7378 27424
rect 7321 26662 7379 26672
rect 7321 26343 7325 26662
rect 7325 26343 7377 26662
rect 7377 26343 7379 26662
rect 7321 26333 7379 26343
rect 3015 25119 3113 25519
rect 4937 25474 5417 25477
rect 4937 25422 5417 25474
rect 4937 25419 5417 25422
rect 7395 25475 7875 25479
rect 7395 25423 7875 25475
rect 7395 25421 7875 25423
rect 12123 27539 12187 28539
rect 13875 27539 13939 28539
rect 12999 26379 13063 27379
rect 15329 29145 15339 29245
rect 15339 29145 15621 29245
rect 21045 27054 21109 27254
rect 23161 27330 23225 27530
rect 25277 27054 25341 27254
rect 27028 27784 27326 28171
rect 21045 26168 21109 26368
rect 23161 25892 23225 26092
rect 25277 26168 25341 26368
rect 9129 23382 9383 23600
rect 12133 24413 12197 24513
rect 19885 24413 19949 24513
rect 16009 24237 16073 24337
rect 16009 24003 16073 24103
rect 12133 23827 12197 23927
rect 19885 23827 19949 23927
rect 11870 23392 11872 23594
rect 11872 23590 12019 23594
rect 12019 23590 19325 23594
rect 11872 23589 12113 23590
rect 12113 23589 19325 23590
rect 11872 23392 19325 23589
rect 11870 23391 19325 23392
rect 19859 23382 20043 23599
rect 16576 22891 16676 23071
rect 16576 22578 16676 22678
rect 11526 20968 11683 21341
rect 12478 21521 12678 21585
rect 13054 21267 13254 21323
rect 13959 20747 14159 20811
rect 12478 19973 12678 20037
rect 13054 20235 13254 20291
rect 14535 21009 14735 21065
rect 14535 20493 14735 20549
rect 13054 19719 13254 19775
rect 13959 19199 14159 19263
rect 12478 18425 12678 18489
rect 13054 18687 13254 18743
rect 14535 19461 14735 19517
rect 14535 18945 14735 19001
rect 13054 18171 13254 18227
rect 13959 17651 14159 17715
rect 12478 16877 12678 16941
rect 13054 17139 13254 17195
rect 14535 17913 14735 17969
rect 14535 17397 14735 17453
rect 13054 16623 13254 16679
rect 13959 16103 14159 16167
rect 13054 15591 13254 15647
rect 14535 16365 14735 16421
rect 14534 15849 14734 15905
rect 12478 15329 12678 15393
rect 16096 18772 16160 18778
rect 16096 18720 16156 18772
rect 16156 18720 16160 18772
rect 16096 18714 16160 18720
rect 23132 24775 23226 24912
rect 22213 24517 22307 24654
rect 24048 24517 24142 24654
rect 20736 24242 20819 24342
rect 20726 24056 20839 24156
rect 22214 23728 22308 23865
rect 24046 23728 24140 23865
rect 21347 23382 21659 23600
rect 23131 23517 23225 23654
rect 24701 22956 24842 23018
rect 29707 24068 29886 24249
rect 22571 22533 22627 22673
rect 20371 18713 20450 18779
rect 30362 20632 30542 20775
rect 18099 17743 18521 18131
rect 30367 17477 30537 17647
rect 16883 16852 17023 16916
rect 15374 16726 15447 16806
rect 16883 16336 17023 16400
rect 15580 15941 16180 16015
rect 16763 15749 16828 16108
rect 16763 15295 16828 15654
rect 30362 12891 30542 13028
rect 13963 11892 14168 12273
rect 1903 10020 2303 10420
rect 3113 10136 3313 10200
rect 3689 9882 3889 9938
rect 4594 9362 4794 9426
rect 3113 8588 3313 8652
rect 3689 8850 3889 8906
rect 5169 9624 5369 9680
rect 5170 9108 5370 9164
rect 3689 8334 3889 8390
rect 4594 7814 4794 7878
rect 3113 7040 3313 7104
rect 3689 7302 3889 7358
rect 5170 8076 5370 8132
rect 5170 7560 5370 7616
rect 3689 6786 3889 6842
rect 4594 6266 4794 6330
rect 3113 5492 3313 5556
rect 3689 5754 3889 5810
rect 5170 6528 5370 6584
rect 5170 6012 5370 6068
rect 3689 5238 3889 5294
rect 4594 4718 4794 4782
rect 3113 3944 3313 4008
rect 3689 4206 3889 4262
rect 5170 4980 5370 5036
rect 5170 4464 5370 4520
rect 6215 9514 6815 9588
rect 7398 9875 7463 10234
rect 7398 9421 7463 9780
rect 7518 9129 7658 9193
rect 5997 8666 6082 8746
rect 7518 8613 7658 8677
rect 25902 11004 26136 11404
rect 18058 7286 18634 7296
rect 18058 7231 18634 7286
rect 11501 6169 11886 6554
rect 18673 6239 18676 7037
rect 18676 6239 18728 7037
rect 18728 6239 18731 7037
rect 26498 9303 26678 9458
rect 21831 7957 21887 7970
rect 21831 7638 21835 7957
rect 21835 7638 21887 7957
rect 21831 7628 21887 7638
rect 30362 8087 30542 8230
rect 21830 6876 21888 6886
rect 21830 6557 21834 6876
rect 21834 6557 21886 6876
rect 21886 6557 21888 6876
rect 21830 6547 21888 6557
rect 19446 5688 19926 5691
rect 19446 5636 19926 5688
rect 19446 5633 19926 5636
rect 21904 5689 22384 5693
rect 21904 5637 22384 5689
rect 21904 5635 22384 5637
rect 7178 2658 7358 2767
<< metal3 >>
rect 11855 32983 14354 32988
rect 11855 32876 11865 32983
rect 14344 32876 14354 32983
rect 11855 32871 14354 32876
rect 12989 31777 13073 31782
rect 10925 31121 11675 31126
rect 10925 30961 10935 31121
rect 11665 30961 11675 31121
rect 10925 30956 11675 30961
rect 12989 30777 12999 31777
rect 13063 30863 13073 31777
rect 16564 31278 18644 31298
rect 16564 31214 16592 31278
rect 18616 31214 18644 31278
rect 13063 30777 14181 30863
rect 12989 30772 14181 30777
rect 13003 30763 14181 30772
rect 12112 30540 12196 30545
rect 12112 29540 12122 30540
rect 12186 29540 12196 30540
rect 12112 29535 12196 29540
rect 13865 30540 13949 30545
rect 13865 29540 13875 30540
rect 13939 29540 13949 30540
rect 13865 29535 13949 29540
rect 14081 28547 14181 30763
rect 16564 29947 18644 31214
rect 16564 29767 26614 29947
rect 16564 29250 18644 29767
rect 15319 29245 18644 29250
rect 15319 29145 15329 29245
rect 15621 29145 18644 29245
rect 15319 29140 18644 29145
rect 16564 28926 18644 29140
rect 14081 28544 14272 28547
rect 12113 28539 14272 28544
rect 7311 27756 7389 27761
rect 7311 27414 7322 27756
rect 7378 27414 7389 27756
rect 12113 27539 12123 28539
rect 12187 28444 13875 28539
rect 12187 27539 12197 28444
rect 12113 27534 12197 27539
rect 13865 27539 13875 28444
rect 13939 28444 14272 28539
rect 13939 27539 13949 28444
rect 13865 27534 13949 27539
rect 7311 27087 7389 27414
rect 3539 27082 7389 27087
rect 3539 27017 3549 27082
rect 4125 27017 7389 27082
rect 3539 27012 7389 27017
rect 4154 26823 4334 26828
rect 4154 26025 4164 26823
rect 4222 26025 4334 26823
rect 7311 26672 7389 27012
rect 7311 26333 7321 26672
rect 7379 26333 7389 26672
rect 12989 27379 13073 27384
rect 12989 26379 12999 27379
rect 13063 26379 13073 27379
rect 12989 26374 13073 26379
rect 7311 26328 7389 26333
rect 3005 25519 3123 25524
rect 3005 25119 3015 25519
rect 3113 25119 3123 25519
rect 3005 25114 3123 25119
rect 4154 25059 4334 26025
rect 4927 25477 5427 25482
rect 4927 25419 4937 25477
rect 5417 25419 5427 25477
rect 4927 25414 5427 25419
rect 7385 25479 7885 25484
rect 7385 25421 7395 25479
rect 7875 25421 7885 25479
rect 7385 25416 7885 25421
rect 4144 24955 4154 25059
rect 4334 24955 4344 25059
rect 4154 24860 4334 24955
rect 4927 12970 5107 25414
rect 7385 13785 7565 25416
rect 12116 24513 12214 24518
rect 12116 24413 12133 24513
rect 12197 24413 12214 24513
rect 12116 24408 12214 24413
rect 14162 24342 14272 28444
rect 23151 27530 23235 27535
rect 23151 27330 23161 27530
rect 23225 27330 23235 27530
rect 23151 27325 23235 27330
rect 21035 27254 21119 27259
rect 21035 27054 21045 27254
rect 21109 27149 21119 27254
rect 25267 27254 25351 27259
rect 25267 27149 25277 27254
rect 21109 27054 25277 27149
rect 25341 27149 25351 27254
rect 25341 27054 25791 27149
rect 21035 27049 25791 27054
rect 21035 26368 21119 26373
rect 21035 26168 21045 26368
rect 21109 26168 21119 26368
rect 21035 26163 21119 26168
rect 25267 26368 25351 26373
rect 25267 26168 25277 26368
rect 25341 26168 25351 26368
rect 25267 26163 25351 26168
rect 23151 26092 23235 26097
rect 23151 25892 23161 26092
rect 23225 25987 23235 26092
rect 25691 25987 25791 27049
rect 23225 25892 25791 25987
rect 23151 25887 25791 25892
rect 23122 24912 23236 24917
rect 23122 24775 23132 24912
rect 23226 24775 23236 24912
rect 23122 24770 23236 24775
rect 24321 24659 24468 25887
rect 22203 24654 24468 24659
rect 19847 24513 19975 24518
rect 19847 24413 19885 24513
rect 19949 24413 19975 24513
rect 22203 24517 22213 24654
rect 22307 24517 24048 24654
rect 24142 24517 24468 24654
rect 22203 24512 24468 24517
rect 19847 24408 19975 24413
rect 20726 24342 20829 24347
rect 14162 24337 20345 24342
rect 14162 24237 16009 24337
rect 16073 24237 20345 24337
rect 20695 24242 20736 24342
rect 20819 24242 20829 24342
rect 20726 24237 20829 24242
rect 14162 24232 20345 24237
rect 20235 24156 20345 24232
rect 20716 24156 20849 24161
rect 15983 24103 16098 24108
rect 15983 24003 16009 24103
rect 16073 24003 16098 24103
rect 15983 23998 16098 24003
rect 20235 24056 20726 24156
rect 20839 24056 20849 24156
rect 20235 23932 20345 24056
rect 20716 24051 20849 24056
rect 12123 23927 20345 23932
rect 12123 23827 12133 23927
rect 12197 23827 19885 23927
rect 19949 23827 20345 23927
rect 12123 23822 20345 23827
rect 22204 23865 22318 23870
rect 22204 23728 22214 23865
rect 22308 23728 22318 23865
rect 22204 23723 22318 23728
rect 24036 23865 24150 23870
rect 24036 23728 24046 23865
rect 24140 23728 24150 23865
rect 24036 23723 24150 23728
rect 23121 23654 23235 23659
rect 24321 23654 24468 24512
rect 9119 23600 9393 23605
rect 9119 23382 9129 23600
rect 9383 23382 9393 23600
rect 19849 23599 20053 23604
rect 11860 23594 19335 23599
rect 11860 23391 11870 23594
rect 19325 23391 19335 23594
rect 11860 23386 19335 23391
rect 9119 23377 9393 23382
rect 19849 23382 19859 23599
rect 20043 23382 20053 23599
rect 19849 23377 20053 23382
rect 21337 23600 21669 23605
rect 21337 23382 21347 23600
rect 21659 23382 21669 23600
rect 23121 23517 23131 23654
rect 23225 23517 24468 23654
rect 23121 23512 24468 23517
rect 21337 23377 21669 23382
rect 16566 23071 16686 23076
rect 16566 22891 16576 23071
rect 16676 22891 16686 23071
rect 24691 23021 24852 23023
rect 24691 22953 24701 23021
rect 24842 22953 24852 23021
rect 24691 22951 24852 22953
rect 16566 22886 16686 22891
rect 16566 22678 16686 22683
rect 16566 22578 16576 22678
rect 16676 22673 22637 22678
rect 16676 22578 22571 22673
rect 16566 22573 16686 22578
rect 22561 22533 22571 22578
rect 22627 22533 22637 22673
rect 22561 22528 22637 22533
rect 26434 22432 26614 29767
rect 27018 28171 27336 28176
rect 27018 27784 27028 28171
rect 27326 27784 27336 28171
rect 27018 27779 27336 27784
rect 29697 24249 29896 24254
rect 29697 24068 29707 24249
rect 29886 24068 29896 24249
rect 29697 24063 29896 24068
rect 24403 22404 28175 22432
rect 12473 21585 12683 21595
rect 12473 21521 12478 21585
rect 12678 21521 12683 21585
rect 12473 21511 12683 21521
rect 24403 21459 28091 22404
rect 24181 21352 28091 21459
rect 11516 21341 11693 21346
rect 11516 20968 11526 21341
rect 11683 20968 11693 21341
rect 13049 21323 13259 21333
rect 13049 21267 13054 21323
rect 13254 21267 13259 21323
rect 13049 21257 13259 21267
rect 11516 20963 11693 20968
rect 13183 21193 13259 21257
rect 13183 20301 13257 21193
rect 14530 21065 14740 21075
rect 14530 21009 14535 21065
rect 14735 21009 14740 21065
rect 14530 20999 14740 21009
rect 13954 20811 14164 20821
rect 13954 20747 13959 20811
rect 14159 20747 14164 20811
rect 13954 20737 14164 20747
rect 14664 20559 14740 20999
rect 14530 20549 14740 20559
rect 14530 20493 14535 20549
rect 14735 20493 14740 20549
rect 14530 20483 14740 20493
rect 13049 20291 13259 20301
rect 13049 20235 13054 20291
rect 13254 20235 13259 20291
rect 13049 20225 13259 20235
rect 12473 20037 12683 20047
rect 12473 19973 12478 20037
rect 12678 19973 12683 20037
rect 12473 19963 12683 19973
rect 13183 19785 13257 20225
rect 13049 19775 13259 19785
rect 13049 19719 13054 19775
rect 13254 19719 13259 19775
rect 13049 19709 13259 19719
rect 13183 18753 13257 19709
rect 14664 19527 14740 20483
rect 14530 19517 14740 19527
rect 14530 19461 14535 19517
rect 14735 19461 14740 19517
rect 14530 19451 14740 19461
rect 13954 19263 14164 19273
rect 13954 19199 13959 19263
rect 14159 19199 14164 19263
rect 13954 19189 14164 19199
rect 14664 19011 14740 19451
rect 14530 19001 14740 19011
rect 14530 18945 14535 19001
rect 14735 18945 14740 19001
rect 24403 18980 28091 21352
rect 28155 18980 28175 22404
rect 30352 20775 30552 20780
rect 30352 20632 30362 20775
rect 30542 20632 30552 20775
rect 30352 20627 30552 20632
rect 24403 18952 28175 18980
rect 14530 18935 14740 18945
rect 13049 18743 13259 18753
rect 13049 18687 13054 18743
rect 13254 18687 13259 18743
rect 13049 18677 13259 18687
rect 12473 18489 12683 18499
rect 12473 18425 12478 18489
rect 12678 18425 12683 18489
rect 12473 18415 12683 18425
rect 13183 18237 13257 18677
rect 13049 18227 13259 18237
rect 13049 18171 13054 18227
rect 13254 18171 13259 18227
rect 13049 18161 13259 18171
rect 13183 17205 13257 18161
rect 14664 17979 14740 18935
rect 16091 18778 16208 18788
rect 16091 18714 16096 18778
rect 16160 18714 16208 18778
rect 16091 18704 16208 18714
rect 20344 18779 20467 18786
rect 20344 18713 20371 18779
rect 20450 18713 20467 18779
rect 20344 18702 20467 18713
rect 14530 17969 14740 17979
rect 14530 17913 14535 17969
rect 14735 17913 14740 17969
rect 14530 17903 14740 17913
rect 13954 17715 14164 17725
rect 13954 17651 13959 17715
rect 14159 17651 14164 17715
rect 13954 17641 14164 17651
rect 14664 17463 14740 17903
rect 18089 18131 18531 18136
rect 18089 17743 18099 18131
rect 18521 17743 18531 18131
rect 18089 17738 18531 17743
rect 30363 17652 30541 17657
rect 30362 17651 30542 17652
rect 30362 17473 30363 17651
rect 30541 17473 30542 17651
rect 30362 17472 30542 17473
rect 30363 17467 30541 17472
rect 14530 17453 14740 17463
rect 14530 17397 14535 17453
rect 14735 17397 14740 17453
rect 14530 17387 14740 17397
rect 13049 17195 13259 17205
rect 13049 17139 13054 17195
rect 13254 17139 13259 17195
rect 13049 17129 13259 17139
rect 12473 16941 12683 16951
rect 12473 16877 12478 16941
rect 12678 16877 12683 16941
rect 12473 16867 12683 16877
rect 13183 16689 13257 17129
rect 13049 16679 13259 16689
rect 13049 16623 13054 16679
rect 13254 16623 13259 16679
rect 13049 16613 13259 16623
rect 13183 15657 13257 16613
rect 14664 16507 14740 17387
rect 16878 16916 17028 16926
rect 16878 16852 16883 16916
rect 17023 16852 17028 16916
rect 16878 16842 17028 16852
rect 15369 16806 15452 16816
rect 15369 16726 15374 16806
rect 15447 16726 15452 16806
rect 15369 16716 15452 16726
rect 15374 16507 15447 16716
rect 14664 16431 15447 16507
rect 14530 16421 14740 16431
rect 14530 16365 14535 16421
rect 14735 16365 14740 16421
rect 14530 16355 14740 16365
rect 13954 16167 14164 16177
rect 13954 16103 13959 16167
rect 14159 16103 14164 16167
rect 13954 16093 14164 16103
rect 14664 15915 14740 16355
rect 16878 16400 17028 16410
rect 16878 16336 16883 16400
rect 17023 16336 17028 16400
rect 16878 16326 17028 16336
rect 16758 16108 16833 16118
rect 15575 16015 16185 16025
rect 15575 15941 15580 16015
rect 16180 15941 16185 16015
rect 15575 15931 16185 15941
rect 14529 15905 14740 15915
rect 14529 15849 14534 15905
rect 14734 15849 14740 15905
rect 14529 15839 14740 15849
rect 13049 15647 13259 15657
rect 13049 15591 13054 15647
rect 13254 15591 13259 15647
rect 13049 15581 13259 15591
rect 12473 15393 12683 15403
rect 12473 15329 12478 15393
rect 12678 15329 12683 15393
rect 12473 15319 12683 15329
rect 13183 15265 13257 15581
rect 14664 15265 14740 15839
rect 16758 15749 16763 16108
rect 16828 15749 16833 16108
rect 16758 15739 16833 15749
rect 16758 15654 16833 15664
rect 16758 15295 16763 15654
rect 16828 15295 16833 15654
rect 16758 15285 16833 15295
rect 13183 15191 14740 15265
rect 7385 13605 11623 13785
rect 11772 13605 11782 13785
rect 30352 13028 30552 13033
rect 4927 12790 9240 12970
rect 9417 12790 9427 12970
rect 30352 12891 30362 13028
rect 30542 12891 30552 13028
rect 30352 12886 30552 12891
rect 13953 12273 14178 12278
rect 13953 11892 13963 12273
rect 14168 11892 14178 12273
rect 13953 11887 14178 11892
rect 4867 11174 4873 11559
rect 5258 11174 11886 11559
rect 1893 10420 2313 10425
rect 1893 10020 1903 10420
rect 2303 10020 2313 10420
rect 3818 10264 5375 10338
rect 3108 10200 3318 10210
rect 3108 10136 3113 10200
rect 3313 10136 3318 10200
rect 3108 10126 3318 10136
rect 1893 10015 2313 10020
rect 3818 9948 3892 10264
rect 3684 9938 3894 9948
rect 3684 9882 3689 9938
rect 3889 9882 3894 9938
rect 3684 9872 3894 9882
rect 3818 8916 3892 9872
rect 5299 9690 5375 10264
rect 7393 10234 7468 10244
rect 7393 9875 7398 10234
rect 7463 9875 7468 10234
rect 7393 9865 7468 9875
rect 5164 9680 5375 9690
rect 5164 9624 5169 9680
rect 5369 9624 5375 9680
rect 5164 9614 5375 9624
rect 4589 9426 4799 9436
rect 4589 9362 4594 9426
rect 4794 9362 4799 9426
rect 4589 9352 4799 9362
rect 5299 9174 5375 9614
rect 7393 9780 7468 9790
rect 6210 9588 6820 9598
rect 6210 9514 6215 9588
rect 6815 9514 6820 9588
rect 6210 9504 6820 9514
rect 7393 9421 7398 9780
rect 7463 9421 7468 9780
rect 7393 9411 7468 9421
rect 5165 9164 5375 9174
rect 5165 9108 5170 9164
rect 5370 9108 5375 9164
rect 7513 9193 7663 9203
rect 7513 9129 7518 9193
rect 7658 9129 7663 9193
rect 7513 9119 7663 9129
rect 5165 9098 5375 9108
rect 5299 9022 6082 9098
rect 3684 8906 3894 8916
rect 3684 8850 3689 8906
rect 3889 8850 3894 8906
rect 3684 8840 3894 8850
rect 3108 8652 3318 8662
rect 3108 8588 3113 8652
rect 3313 8588 3318 8652
rect 3108 8578 3318 8588
rect 3818 8400 3892 8840
rect 3684 8390 3894 8400
rect 3684 8334 3689 8390
rect 3889 8334 3894 8390
rect 3684 8324 3894 8334
rect 3818 7368 3892 8324
rect 5299 8142 5375 9022
rect 5997 8756 6082 9022
rect 5992 8746 6087 8756
rect 5992 8666 5997 8746
rect 6082 8666 6087 8746
rect 5992 8656 6087 8666
rect 7513 8677 7663 8687
rect 7513 8613 7518 8677
rect 7658 8613 7663 8677
rect 7513 8603 7663 8613
rect 5165 8132 5375 8142
rect 5165 8076 5170 8132
rect 5370 8076 5375 8132
rect 5165 8066 5375 8076
rect 4589 7878 4799 7888
rect 4589 7814 4594 7878
rect 4794 7814 4799 7878
rect 4589 7804 4799 7814
rect 5299 7626 5375 8066
rect 5165 7616 5375 7626
rect 5165 7560 5170 7616
rect 5370 7560 5375 7616
rect 5165 7550 5375 7560
rect 3684 7358 3894 7368
rect 3684 7302 3689 7358
rect 3889 7302 3894 7358
rect 3684 7292 3894 7302
rect 3108 7104 3318 7114
rect 3108 7040 3113 7104
rect 3313 7040 3318 7104
rect 3108 7030 3318 7040
rect 3818 6852 3892 7292
rect 3684 6842 3894 6852
rect 3684 6786 3689 6842
rect 3889 6786 3894 6842
rect 3684 6776 3894 6786
rect 3818 5820 3892 6776
rect 5299 6594 5375 7550
rect 5165 6584 5375 6594
rect 5165 6528 5170 6584
rect 5370 6528 5375 6584
rect 11501 6559 11886 11174
rect 25892 11404 26146 11409
rect 25892 11004 25902 11404
rect 26136 11004 26146 11404
rect 25892 10999 26146 11004
rect 26488 9458 26688 9463
rect 26488 9303 26498 9458
rect 26678 9303 26688 9458
rect 26488 9298 26688 9303
rect 30352 8230 30552 8235
rect 30352 8087 30362 8230
rect 30542 8087 30552 8230
rect 30352 8082 30552 8087
rect 21820 7970 21898 7975
rect 21820 7628 21831 7970
rect 21887 7628 21898 7970
rect 21820 7301 21898 7628
rect 18048 7296 21898 7301
rect 18048 7231 18058 7296
rect 18634 7231 21898 7296
rect 18048 7226 21898 7231
rect 18663 7037 18843 7042
rect 5165 6518 5375 6528
rect 4589 6330 4799 6340
rect 4589 6266 4594 6330
rect 4794 6266 4799 6330
rect 4589 6256 4799 6266
rect 5299 6078 5375 6518
rect 11496 6554 11891 6559
rect 11496 6169 11501 6554
rect 11886 6169 11891 6554
rect 11496 6164 11891 6169
rect 18663 6239 18673 7037
rect 18731 6239 18843 7037
rect 21820 6886 21898 7226
rect 21820 6547 21830 6886
rect 21888 6547 21898 6886
rect 21820 6542 21898 6547
rect 5165 6068 5375 6078
rect 5165 6012 5170 6068
rect 5370 6012 5375 6068
rect 5165 6002 5375 6012
rect 3684 5810 3894 5820
rect 3684 5754 3689 5810
rect 3889 5754 3894 5810
rect 3684 5744 3894 5754
rect 3108 5556 3318 5566
rect 3108 5492 3113 5556
rect 3313 5492 3318 5556
rect 3108 5482 3318 5492
rect 3818 5304 3892 5744
rect 3684 5294 3894 5304
rect 3684 5238 3689 5294
rect 3889 5238 3894 5294
rect 3684 5228 3894 5238
rect 3818 4336 3892 5228
rect 5299 5046 5375 6002
rect 5165 5036 5375 5046
rect 5165 4980 5170 5036
rect 5370 4980 5375 5036
rect 5165 4970 5375 4980
rect 4589 4782 4799 4792
rect 4589 4718 4594 4782
rect 4794 4718 4799 4782
rect 4589 4708 4799 4718
rect 5299 4530 5375 4970
rect 5165 4520 5375 4530
rect 5165 4464 5170 4520
rect 5370 4464 5375 4520
rect 5165 4454 5375 4464
rect 3818 4272 3894 4336
rect 3684 4262 3894 4272
rect 3684 4206 3689 4262
rect 3889 4206 3894 4262
rect 3684 4196 3894 4206
rect 3108 4008 3318 4018
rect 3108 3944 3113 4008
rect 3313 3944 3318 4008
rect 3108 3934 3318 3944
rect 18663 3571 18843 6239
rect 14906 3391 18843 3571
rect 19436 5691 19936 5696
rect 19436 5633 19446 5691
rect 19926 5633 19936 5691
rect 19436 5628 19936 5633
rect 21894 5693 22394 5698
rect 21894 5635 21904 5693
rect 22384 5635 22394 5693
rect 21894 5630 22394 5635
rect 7168 2767 7368 2772
rect 7168 2658 7178 2767
rect 7358 2658 7368 2767
rect 7168 2653 7368 2658
rect 14906 1818 15086 3391
rect 19436 2805 19616 5628
rect 21894 4301 22074 5630
rect 21884 4121 21894 4301
rect 22074 4121 22084 4301
rect 21894 4119 22074 4121
rect 19426 2625 19436 2805
rect 19616 2625 19626 2805
rect 14896 1638 14906 1818
rect 15086 1638 15096 1818
<< via3 >>
rect 11865 32876 14344 32983
rect 10935 30961 11665 31121
rect 16592 31214 18616 31278
rect 12122 29540 12186 30540
rect 13875 29540 13939 30540
rect 12999 26379 13063 27379
rect 3015 25119 3113 25519
rect 4154 24955 4334 25059
rect 12133 24413 12197 24513
rect 23161 27330 23225 27530
rect 21045 26168 21109 26368
rect 25277 26168 25341 26368
rect 23132 24775 23226 24912
rect 19885 24413 19949 24513
rect 20736 24242 20819 24342
rect 16009 24003 16073 24103
rect 20726 24056 20839 24156
rect 22214 23728 22308 23865
rect 24046 23728 24140 23865
rect 9129 23382 9383 23600
rect 11870 23391 19325 23594
rect 19859 23382 20043 23599
rect 21347 23382 21659 23600
rect 16576 22891 16676 23071
rect 24701 23018 24842 23021
rect 24701 22956 24842 23018
rect 24701 22953 24842 22956
rect 27028 27784 27326 28171
rect 29707 24068 29886 24249
rect 12478 21521 12678 21585
rect 11526 20968 11683 21341
rect 13959 20747 14159 20811
rect 12478 19973 12678 20037
rect 13959 19199 14159 19263
rect 28091 18980 28155 22404
rect 30362 20632 30542 20775
rect 12478 18425 12678 18489
rect 16096 18714 16160 18778
rect 20371 18713 20450 18779
rect 13959 17651 14159 17715
rect 18099 17743 18521 18131
rect 30363 17647 30541 17651
rect 30363 17477 30367 17647
rect 30367 17477 30537 17647
rect 30537 17477 30541 17647
rect 30363 17473 30541 17477
rect 12478 16877 12678 16941
rect 16883 16852 17023 16916
rect 13959 16103 14159 16167
rect 16883 16336 17023 16400
rect 15580 15941 16180 16015
rect 12478 15329 12678 15393
rect 16763 15749 16828 16108
rect 16763 15295 16828 15654
rect 11623 13605 11772 13785
rect 9240 12790 9417 12970
rect 30362 12891 30542 13028
rect 13963 11892 14168 12273
rect 4873 11174 5258 11559
rect 1903 10020 2303 10420
rect 3113 10136 3313 10200
rect 7398 9875 7463 10234
rect 4594 9362 4794 9426
rect 6215 9514 6815 9588
rect 7398 9421 7463 9780
rect 7518 9129 7658 9193
rect 3113 8588 3313 8652
rect 7518 8613 7658 8677
rect 4594 7814 4794 7878
rect 3113 7040 3313 7104
rect 25902 11004 26136 11404
rect 26498 9303 26678 9458
rect 30362 8087 30542 8230
rect 4594 6266 4794 6330
rect 3113 5492 3313 5556
rect 4594 4718 4794 4782
rect 3113 3944 3313 4008
rect 7178 2658 7358 2767
rect 21894 4121 22074 4301
rect 19436 2625 19616 2805
rect 14906 1638 15086 1818
<< mimcap >>
rect 16604 30926 18604 30966
rect 16604 29006 16644 30926
rect 18564 29006 18604 30926
rect 16604 28966 18604 29006
rect 24443 22352 27843 22392
rect 24443 19032 24483 22352
rect 27803 19032 27843 22352
rect 24443 18992 27843 19032
<< mimcapcontact >>
rect 16644 29006 18564 30926
rect 24483 19032 27803 22352
<< metal4 >>
rect 400 43919 800 44152
rect 400 43282 2000 43919
rect 400 25519 800 43282
rect 31400 33199 31800 44152
rect 14344 33198 31800 33199
rect 11711 33197 31800 33198
rect 11470 32983 31800 33197
rect 11470 32876 11865 32983
rect 14344 32876 31800 32983
rect 11470 32798 31800 32876
rect 11470 31122 11930 32798
rect 14502 32797 31800 32798
rect 16576 31278 18632 31294
rect 16576 31214 16592 31278
rect 18616 31214 18632 31278
rect 16576 31198 18632 31214
rect 10934 31121 11930 31122
rect 10934 30961 10935 31121
rect 11665 30961 11930 31121
rect 10934 30960 11930 30961
rect 11470 30794 11930 30960
rect 16643 30926 18565 30927
rect 12121 30540 12187 30541
rect 12121 29540 12122 30540
rect 12186 29639 12187 30540
rect 13874 30540 13940 30541
rect 13874 29639 13875 30540
rect 12186 29540 13875 29639
rect 13939 29639 13940 30540
rect 13939 29540 14575 29639
rect 12121 29539 14575 29540
rect 12998 27379 13064 27380
rect 12998 26379 12999 27379
rect 13063 27345 13064 27379
rect 14475 27345 14575 29539
rect 16643 29006 16644 30926
rect 18564 29110 18565 30926
rect 31400 30560 31800 32797
rect 31399 30160 31800 30560
rect 18564 29044 19967 29110
rect 18564 29006 18565 29044
rect 16643 29005 18565 29006
rect 13063 27245 14575 27345
rect 19901 27331 19967 29044
rect 31400 28175 31800 30160
rect 27027 28171 27327 28172
rect 29046 28171 31800 28175
rect 26765 27784 27028 28171
rect 27326 27784 31800 28171
rect 27027 27783 27327 27784
rect 28887 27621 31800 27784
rect 13063 26379 13064 27245
rect 12998 26378 13064 26379
rect 3014 25519 3114 25520
rect 400 25119 3015 25519
rect 3113 25119 3189 25519
rect 400 23600 800 25119
rect 3014 25118 3114 25119
rect 4153 25059 4335 25060
rect 4153 24955 4154 25059
rect 4334 24955 4335 25059
rect 4153 24954 4335 24955
rect 4154 24837 4334 24954
rect 4154 24657 10288 24837
rect 9128 23600 9384 23601
rect 400 23382 9129 23600
rect 9383 23382 9384 23600
rect 400 11559 800 23382
rect 8157 21341 8530 23382
rect 9128 23381 9384 23382
rect 10108 23071 10288 24657
rect 14475 24514 14575 27245
rect 19900 27253 19967 27331
rect 20592 27530 23226 27531
rect 20592 27431 23161 27530
rect 19900 24514 19966 27253
rect 20592 26369 20692 27431
rect 23160 27330 23161 27431
rect 23225 27330 23226 27530
rect 23160 27329 23226 27330
rect 20592 26368 25342 26369
rect 20592 26269 21045 26368
rect 21044 26168 21045 26269
rect 21109 26269 25277 26368
rect 21109 26168 21110 26269
rect 21044 26167 21110 26168
rect 21937 24913 22076 26269
rect 25276 26168 25277 26269
rect 25341 26168 25342 26368
rect 25276 26167 25342 26168
rect 21937 24912 23249 24913
rect 21937 24775 23132 24912
rect 23226 24775 23249 24912
rect 21937 24774 23249 24775
rect 12132 24513 20613 24514
rect 12132 24413 12133 24513
rect 12197 24413 19885 24513
rect 19949 24413 20613 24513
rect 12132 24412 20613 24413
rect 20511 24342 20613 24412
rect 20735 24342 20820 24343
rect 20511 24242 20736 24342
rect 20819 24242 20820 24342
rect 20511 24104 20613 24242
rect 20735 24241 20820 24242
rect 20725 24156 20840 24157
rect 16008 24103 20613 24104
rect 16008 24003 16009 24103
rect 16073 24003 20613 24103
rect 20701 24056 20726 24156
rect 20839 24056 20840 24156
rect 20725 24055 20840 24056
rect 16008 24002 20613 24003
rect 21937 23866 22076 24774
rect 21937 23865 24141 23866
rect 21937 23728 22214 23865
rect 22308 23728 24046 23865
rect 24140 23728 24141 23865
rect 21937 23727 24141 23728
rect 21346 23600 21660 23601
rect 19288 23599 21347 23600
rect 19288 23595 19859 23599
rect 11869 23594 19859 23595
rect 11869 23391 11870 23594
rect 19325 23391 19859 23594
rect 11869 23390 19859 23391
rect 19288 23384 19859 23390
rect 19673 23382 19859 23384
rect 20043 23382 21347 23599
rect 21659 23382 22131 23600
rect 19858 23381 20044 23382
rect 21346 23381 21660 23382
rect 16575 23071 16677 23072
rect 10108 22891 16576 23071
rect 16676 22891 16687 23071
rect 24692 23021 24843 23022
rect 24692 22953 24701 23021
rect 24842 23018 24843 23021
rect 24842 22956 24911 23018
rect 24842 22953 24843 22956
rect 24692 22952 24843 22953
rect 16575 22890 16677 22891
rect 24692 22353 24803 22952
rect 28075 22404 28171 22420
rect 24482 22352 27804 22353
rect 12477 21585 12679 21586
rect 12477 21521 12478 21585
rect 12678 21521 12679 21585
rect 12477 21520 12679 21521
rect 11525 21341 11684 21342
rect 8157 20968 11526 21341
rect 11683 20968 11684 21341
rect 11525 20967 11684 20968
rect 12477 20038 12553 21520
rect 13958 20811 14160 20812
rect 13958 20747 13959 20811
rect 14159 20747 14160 20811
rect 13958 20746 14160 20747
rect 12477 20037 12679 20038
rect 12477 19973 12478 20037
rect 12678 19973 12679 20037
rect 12477 19972 12679 19973
rect 12477 18490 12553 19972
rect 13958 19264 14034 20746
rect 13958 19263 14160 19264
rect 13958 19199 13959 19263
rect 14159 19199 14160 19263
rect 13958 19198 14160 19199
rect 12477 18489 12679 18490
rect 12477 18425 12478 18489
rect 12678 18425 12679 18489
rect 12477 18424 12679 18425
rect 12477 16942 12553 18424
rect 13958 17716 14034 19198
rect 24482 19032 24483 22352
rect 27803 19032 27804 22352
rect 24482 19031 27804 19032
rect 28075 18980 28091 22404
rect 28155 18980 28171 22404
rect 28075 18964 28171 18980
rect 28887 19044 29274 27621
rect 29706 24249 29887 24250
rect 29706 24068 29707 24249
rect 29886 24069 30542 24249
rect 29886 24068 29887 24069
rect 29706 24067 29887 24068
rect 30362 20776 30542 24069
rect 30361 20775 30543 20776
rect 30361 20632 30362 20775
rect 30542 20632 30543 20775
rect 30361 20631 30543 20632
rect 31400 19852 31800 27621
rect 31401 19365 31800 19852
rect 31400 19044 31800 19365
rect 20370 18779 20451 18780
rect 16095 18778 20371 18779
rect 16095 18714 16096 18778
rect 16160 18714 20371 18778
rect 16095 18713 20371 18714
rect 20450 18713 20451 18779
rect 20370 18712 20451 18713
rect 28887 18490 31800 19044
rect 18098 18131 18522 18132
rect 28887 18131 29274 18490
rect 18098 17743 18099 18131
rect 18521 17744 29274 18131
rect 18521 17743 18522 17744
rect 18098 17742 18522 17743
rect 13958 17715 14160 17716
rect 13958 17651 13959 17715
rect 14159 17651 14160 17715
rect 13958 17650 14160 17651
rect 30362 17651 30542 17652
rect 12477 16941 12679 16942
rect 12477 16877 12478 16941
rect 12678 16877 12679 16941
rect 12477 16876 12679 16877
rect 12477 15394 12553 16876
rect 13958 16168 14034 17650
rect 30362 17473 30363 17651
rect 30541 17473 30542 17651
rect 16577 16916 17024 16917
rect 16577 16852 16883 16916
rect 17023 16852 17024 16916
rect 16577 16851 17024 16852
rect 16577 16662 16653 16851
rect 16109 16596 16653 16662
rect 13958 16167 14160 16168
rect 13958 16103 13959 16167
rect 14159 16103 14160 16167
rect 13958 16102 14160 16103
rect 12477 15393 12679 15394
rect 12477 15329 12478 15393
rect 12678 15329 12679 15393
rect 12477 15328 12679 15329
rect 12477 15121 12553 15328
rect 13958 15121 14034 16102
rect 16109 16016 16185 16596
rect 16577 16401 16653 16596
rect 16577 16400 17024 16401
rect 16577 16336 16883 16400
rect 17023 16336 17024 16400
rect 16577 16335 17024 16336
rect 15579 16015 16185 16016
rect 15579 15941 15580 16015
rect 16180 15941 16185 16015
rect 15579 15940 16185 15941
rect 16758 16108 16831 16146
rect 12477 15045 14034 15121
rect 16758 15749 16763 16108
rect 16828 15749 16831 16108
rect 16758 15654 16831 15749
rect 16758 15295 16763 15654
rect 16828 15295 16831 15654
rect 13208 14933 13285 15045
rect 16758 14933 16831 15295
rect 13208 14857 16831 14933
rect 11622 13785 11773 13786
rect 11622 13605 11623 13785
rect 11772 13605 13005 13785
rect 11622 13604 11773 13605
rect 9239 12970 9418 12971
rect 9239 12790 9240 12970
rect 9417 12790 10547 12970
rect 9239 12789 9418 12790
rect 4872 11559 5259 11560
rect 400 11174 4873 11559
rect 5258 11174 5259 11559
rect 400 10420 800 11174
rect 4872 11173 5259 11174
rect 3843 10596 7466 10672
rect 3843 10484 3920 10596
rect 1902 10420 2304 10421
rect 400 10020 1903 10420
rect 2303 10020 2304 10420
rect 400 1000 800 10020
rect 1902 10019 2304 10020
rect 3112 10408 4669 10484
rect 3112 10201 3188 10408
rect 3112 10200 3314 10201
rect 3112 10136 3113 10200
rect 3313 10136 3314 10200
rect 3112 10135 3314 10136
rect 3112 8653 3188 10135
rect 4593 9427 4669 10408
rect 7393 10234 7466 10596
rect 7393 9875 7398 10234
rect 7463 9875 7466 10234
rect 7393 9780 7466 9875
rect 6214 9588 6820 9589
rect 6214 9514 6215 9588
rect 6815 9514 6820 9588
rect 6214 9513 6820 9514
rect 4593 9426 4795 9427
rect 4593 9362 4594 9426
rect 4794 9362 4795 9426
rect 4593 9361 4795 9362
rect 3112 8652 3314 8653
rect 3112 8588 3113 8652
rect 3313 8588 3314 8652
rect 3112 8587 3314 8588
rect 3112 7105 3188 8587
rect 4593 7879 4669 9361
rect 6744 8933 6820 9513
rect 7393 9421 7398 9780
rect 7463 9421 7466 9780
rect 7393 9383 7466 9421
rect 7212 9193 7659 9194
rect 7212 9129 7518 9193
rect 7658 9129 7659 9193
rect 7212 9128 7659 9129
rect 7212 8933 7288 9128
rect 6744 8867 7288 8933
rect 7212 8678 7288 8867
rect 7212 8677 7659 8678
rect 7212 8613 7518 8677
rect 7658 8613 7659 8677
rect 7212 8612 7659 8613
rect 4593 7878 4795 7879
rect 4593 7814 4594 7878
rect 4794 7814 4795 7878
rect 4593 7813 4795 7814
rect 3112 7104 3314 7105
rect 3112 7040 3113 7104
rect 3313 7040 3314 7104
rect 3112 7039 3314 7040
rect 3112 5557 3188 7039
rect 4593 6331 4669 7813
rect 4593 6330 4795 6331
rect 4593 6266 4594 6330
rect 4794 6266 4795 6330
rect 4593 6265 4795 6266
rect 3112 5556 3314 5557
rect 3112 5492 3113 5556
rect 3313 5492 3314 5556
rect 3112 5491 3314 5492
rect 3112 4009 3188 5491
rect 4593 4783 4669 6265
rect 4593 4782 4795 4783
rect 4593 4718 4594 4782
rect 4794 4718 4795 4782
rect 4593 4717 4795 4718
rect 3112 4008 3314 4009
rect 3112 3944 3113 4008
rect 3313 3944 3314 4008
rect 3112 3943 3314 3944
rect 10367 2805 10547 12790
rect 12825 4301 13005 13605
rect 30362 13029 30542 17473
rect 30361 13028 30543 13029
rect 30361 12891 30362 13028
rect 30542 12891 30543 13028
rect 30361 12890 30543 12891
rect 13962 12273 14169 12274
rect 13962 11892 13963 12273
rect 14168 11892 27933 12273
rect 13962 11891 14169 11892
rect 25901 11404 26137 11405
rect 27552 11404 27933 11892
rect 31400 11404 31800 18490
rect 25901 11004 25902 11404
rect 26136 11004 31800 11404
rect 25901 11003 26137 11004
rect 26497 9458 26679 9459
rect 26497 9303 26498 9458
rect 26678 9303 26679 9458
rect 26497 9302 26679 9303
rect 21893 4301 22075 4302
rect 12825 4121 21894 4301
rect 22074 4121 22814 4301
rect 21893 4120 22075 4121
rect 19435 2805 19617 2806
rect 7177 2767 7359 2768
rect 7177 2658 7178 2767
rect 7358 2658 7359 2767
rect 7177 2657 7359 2658
rect 7178 1683 7358 2657
rect 10367 2625 19436 2805
rect 19616 2625 19617 2805
rect 14905 1818 15087 1819
rect 7178 1503 11222 1683
rect 14905 1638 14906 1818
rect 15086 1638 15087 1818
rect 14905 1637 15087 1638
rect 11042 338 11222 1503
rect 11041 199 11222 338
rect 11042 0 11222 199
rect 14906 0 15086 1637
rect 18770 0 18950 2625
rect 19435 2624 19617 2625
rect 22634 0 22814 4121
rect 26498 0 26678 9302
rect 30361 8230 30543 8231
rect 30361 8087 30362 8230
rect 30542 8087 30543 8230
rect 30361 8086 30543 8087
rect 30362 0 30542 8086
rect 31400 1000 31800 11004
<< labels >>
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 31401 1000 31800 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 1000 800 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel metal2 27799 24158 27799 24158 3 3_OTA_0.vo3
rlabel metal3 7464 24429 7464 24429 5 3_OTA_0.vin_p
rlabel metal3 5022 24396 5022 24396 5 3_OTA_0.vin_n
rlabel metal4 14509 33058 14509 33058 3 3_OTA_0.vcc
rlabel metal4 2922 25307 2922 25307 7 3_OTA_0.vss
rlabel metal2 17505 14979 17505 14979 5 3_OTA_0.OTA_vref_0.vcc
rlabel metal2 12146 15011 12146 15011 5 3_OTA_0.OTA_vref_0.vss
rlabel metal2 16619 22612 16619 22612 1 3_OTA_0.OTA_vref_0.vb
rlabel metal4 17695 18747 17695 18747 3 3_OTA_0.OTA_vref_0.vb1
rlabel metal2 17401 17442 17401 17442 1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vcc
rlabel metal2 15810 16968 15810 16968 1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vss
rlabel metal2 16130 16937 16130 16937 1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vref0
rlabel metal1 16810 17370 16810 17370 1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vr
rlabel metal2 16619 22608 16619 22608 1 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vb
rlabel metal4 17687 18743 17687 18743 3 3_OTA_0.OTA_vref_0.OTA_vref_stage2_0.vb1
rlabel metal2 17504 14993 17504 14993 5 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.vcc
rlabel metal2 12140 15021 12140 15021 5 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.vss
rlabel metal3 15444 16464 15444 16464 3 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.vref0
rlabel metal1 16806 17057 16806 17057 1 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.vr
flabel locali 15820 15632 15924 15880 0 FreeSans 400 0 0 0 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter
flabel locali 15249 15691 15298 15792 0 FreeSans 400 0 0 0 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Collector
flabel locali 15408 15668 15448 15786 0 FreeSans 400 0 0 0 3_OTA_0.OTA_vref_0.OTA_vref_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Base
rlabel metal3 7469 24985 7469 24985 5 3_OTA_0.OTA_stage1_0.vin_p
rlabel metal3 5003 24981 5003 24981 5 3_OTA_0.OTA_stage1_0.vin_n
rlabel metal3 4236 24979 4236 24979 5 3_OTA_0.OTA_stage1_0.vb
rlabel metal2 3218 31013 3218 31013 7 3_OTA_0.OTA_stage1_0.vcc
rlabel metal2 3216 25277 3216 25277 7 3_OTA_0.OTA_stage1_0.vss
rlabel metal1 11391 29198 11391 29198 3 3_OTA_0.OTA_stage1_0.vd1
rlabel metal1 11392 28886 11392 28886 3 3_OTA_0.OTA_stage1_0.vd2
rlabel metal2 25778 27996 25778 27996 3 3_OTA_0.3rd_3_OTA_0.vcc
rlabel metal2 22026 21742 22026 21742 7 3_OTA_0.3rd_3_OTA_0.vss
rlabel metal2 26341 24172 26341 24172 3 3_OTA_0.3rd_3_OTA_0.vo3
rlabel metal1 21497 24110 21497 24110 7 3_OTA_0.3rd_3_OTA_0.vd3
rlabel metal1 21497 24287 21497 24287 7 3_OTA_0.3rd_3_OTA_0.vd4
rlabel metal3 24182 21411 24182 21411 7 3_OTA_0.3rd_3_OTA_0.vd1
rlabel metal3 21784 22649 21784 22649 7 3_OTA_0.3rd_3_OTA_0.vb
rlabel metal2 11712 32911 11712 32911 7 3_OTA_0.2nd_3_OTA_0.vcc
rlabel metal2 11808 23485 11808 23485 7 3_OTA_0.2nd_3_OTA_0.vss
rlabel metal1 11607 29197 11607 29197 7 3_OTA_0.2nd_3_OTA_0.vd1
rlabel metal1 11606 28882 11606 28882 7 3_OTA_0.2nd_3_OTA_0.vd2
rlabel metal4 20762 24293 20762 24293 7 3_OTA_0.2nd_3_OTA_0.vd4
rlabel metal3 20761 24105 20761 24105 7 3_OTA_0.2nd_3_OTA_0.vd3
rlabel metal2 20407 23430 20407 23430 5 3_OTA_0.2nd_3_OTA_0.vb1
rlabel metal1 25900 9412 25900 9412 3 diff_final_v0_0.vout
rlabel metal3 21978 5199 21978 5199 5 diff_final_v0_0.vin_p
rlabel metal3 19512 5195 19512 5195 5 diff_final_v0_0.vin_n
rlabel metal3 18745 5193 18745 5193 5 diff_final_v0_0.vb
rlabel metal2 17727 11227 17727 11227 7 diff_final_v0_0.vcc
rlabel metal2 17725 5491 17725 5491 7 diff_final_v0_0.vss
rlabel metal2 7252 2801 7252 2801 1 BGR_BJT_vref_0.vref
rlabel metal2 8141 10572 8141 10572 1 BGR_BJT_vref_0.vcc
rlabel metal2 2775 10558 2775 10558 1 BGR_BJT_vref_0.vss
rlabel metal2 8036 7988 8036 7988 5 BGR_BJT_vref_0.BGR_BJT_stage2_0.vcc
rlabel metal2 6445 8462 6445 8462 5 BGR_BJT_vref_0.BGR_BJT_stage2_0.vss
rlabel metal2 6765 8493 6765 8493 5 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref0
rlabel metal1 7445 8060 7445 8060 5 BGR_BJT_vref_0.BGR_BJT_stage2_0.vr
rlabel metal2 7255 2821 7255 2821 1 BGR_BJT_vref_0.BGR_BJT_stage2_0.vref
rlabel metal2 8139 10536 8139 10536 1 BGR_BJT_vref_0.BGR_BJT_stage1_0.vcc
rlabel metal2 2775 10508 2775 10508 1 BGR_BJT_vref_0.BGR_BJT_stage1_0.vss
rlabel metal3 6079 9065 6079 9065 3 BGR_BJT_vref_0.BGR_BJT_stage1_0.vref0
rlabel metal1 7441 8472 7441 8472 5 BGR_BJT_vref_0.BGR_BJT_stage1_0.vr
flabel locali 6455 9649 6559 9897 0 FreeSans 400 0 0 0 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Emitter
flabel locali 5884 9737 5933 9838 0 FreeSans 400 0 0 0 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Collector
flabel locali 6043 9743 6083 9861 0 FreeSans 400 0 0 0 BGR_BJT_vref_0.BGR_BJT_stage1_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0.Base
<< end >>
